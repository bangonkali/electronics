`timescale 1ns/1ps
module FEAT_INFO_RECT2_ROM(
  addr,
  clk,
  din,
  dout,
  we);

input [11 : 0] addr;
input clk;
input [22 : 0] din;
output reg [22 : 0] dout;
input we;

reg [22:0] mem [0:4095];

initial begin
mem[0]=23'b00000000000000000000000;
mem[1]=23'b00000000000000000000000;
mem[2]=23'b00000000000000000000000;
mem[3]=23'b00000000000000000000000;
mem[4]=23'b00000000000000000000000;
mem[5]=23'b00000000000000000000000;
mem[6]=23'b00000000000000000000000;
mem[7]=23'b00000000000000000000000;
mem[8]=23'b00000000000000000000000;
mem[9]=23'b00000000000000000000000;
mem[10]=23'b00000000000000000000000;
mem[11]=23'b00000000000000000000000;
mem[12]=23'b00000000000000000000000;
mem[13]=23'b00000000000000000000000;
mem[14]=23'b00000000000000000000000;
mem[15]=23'b01000110000100011000110;
mem[16]=23'b00000000000000000000000;
mem[17]=23'b00000000000000000000000;
mem[18]=23'b00000000000000000000000;
mem[19]=23'b00000000000000000000000;
mem[20]=23'b00000000000000000000000;
mem[21]=23'b00000000000000000000000;
mem[22]=23'b00000000000000000000000;
mem[23]=23'b00000000000000000000000;
mem[24]=23'b00000000000000000000000;
mem[25]=23'b00000000000000000000000;
mem[26]=23'b00000000000000000000000;
mem[27]=23'b00000000000000000000000;
mem[28]=23'b00000000000000000000000;
mem[29]=23'b00000000000000000000000;
mem[30]=23'b00000000000000000000000;
mem[31]=23'b01000100010010100101001;
mem[32]=23'b01000010001011000101000;
mem[33]=23'b01000100000100010100101;
mem[34]=23'b01000101001110101100011;
mem[35]=23'b00000000000000000000000;
mem[36]=23'b00000000000000000000000;
mem[37]=23'b00000000000000000000000;
mem[38]=23'b00000000000000000000000;
mem[39]=23'b00000000000000000000000;
mem[40]=23'b00000000000000000000000;
mem[41]=23'b00000000000000000000000;
mem[42]=23'b00000000000000000000000;
mem[43]=23'b00000000000000000000000;
mem[44]=23'b00000000000000000000000;
mem[45]=23'b01000011001000011001011;
mem[46]=23'b00000000000000000000000;
mem[47]=23'b00000000000000000000000;
mem[48]=23'b00000000000000000000000;
mem[49]=23'b01000010001011000101000;
mem[50]=23'b00000000000000000000000;
mem[51]=23'b00000000000000000000000;
mem[52]=23'b00000000000000000000000;
mem[53]=23'b01000101001100100100100;
mem[54]=23'b00000000000000000000000;
mem[55]=23'b00000000000000000000000;
mem[56]=23'b00000000000000000000000;
mem[57]=23'b00000000000000000000000;
mem[58]=23'b01000010000111000100110;
mem[59]=23'b00000000000000000000000;
mem[60]=23'b00000000000000000000000;
mem[61]=23'b00000000000000000000000;
mem[62]=23'b00000000000000000000000;
mem[63]=23'b00000000000000000000000;
mem[64]=23'b00000000000000000000000;
mem[65]=23'b00000000000000000000000;
mem[66]=23'b00000000000000000000000;
mem[67]=23'b00000000000000000000000;
mem[68]=23'b00000000000000000000000;
mem[69]=23'b00000000000000000000000;
mem[70]=23'b00000000000000000000000;
mem[71]=23'b00000000000000000000000;
mem[72]=23'b00000000000000000000000;
mem[73]=23'b00000000000000000000000;
mem[74]=23'b00000000000000000000000;
mem[75]=23'b01000010010010110000001;
mem[76]=23'b00000000000000000000000;
mem[77]=23'b00000000000000000000000;
mem[78]=23'b00000000000000000000000;
mem[79]=23'b00000000000000000000000;
mem[80]=23'b00000000000000000000000;
mem[81]=23'b00000000000000000000000;
mem[82]=23'b00000000000000000000000;
mem[83]=23'b00000000000000000000000;
mem[84]=23'b00000000000000000000000;
mem[85]=23'b00000000000000000000000;
mem[86]=23'b00000000000000000000000;
mem[87]=23'b00000000000000000000000;
mem[88]=23'b00000000000000000000000;
mem[89]=23'b00000000000000000000000;
mem[90]=23'b00000000000000000000000;
mem[91]=23'b00000000000000000000000;
mem[92]=23'b01000010000100001001001;
mem[93]=23'b00000000000000000000000;
mem[94]=23'b00000000000000000000000;
mem[95]=23'b00000000000000000000000;
mem[96]=23'b00000000000000000000000;
mem[97]=23'b00000000000000000000000;
mem[98]=23'b00000000000000000000000;
mem[99]=23'b00000000000000000000000;
mem[100]=23'b00000000000000000000000;
mem[101]=23'b00000000000000000000000;
mem[102]=23'b00000000000000000000000;
mem[103]=23'b00000000000000000000000;
mem[104]=23'b00000000000000000000000;
mem[105]=23'b00000000000000000000000;
mem[106]=23'b01000010000100001001000;
mem[107]=23'b00000000000000000000000;
mem[108]=23'b00000000000000000000000;
mem[109]=23'b01000110001010101001010;
mem[110]=23'b00000000000000000000000;
mem[111]=23'b01000111001100100101000;
mem[112]=23'b00000000000000000000000;
mem[113]=23'b00000000000000000000000;
mem[114]=23'b00000000000000000000000;
mem[115]=23'b00000000000000000000000;
mem[116]=23'b00000000000000000000000;
mem[117]=23'b00000000000000000000000;
mem[118]=23'b01000101000110011100110;
mem[119]=23'b00000000000000000000000;
mem[120]=23'b01000011001001000100111;
mem[121]=23'b00000000000000000000000;
mem[122]=23'b00000000000000000000000;
mem[123]=23'b00000000000000000000000;
mem[124]=23'b01000011001110110001001;
mem[125]=23'b00000000000000000000000;
mem[126]=23'b01000100001000110101010;
mem[127]=23'b00000000000000000000000;
mem[128]=23'b00000000000000000000000;
mem[129]=23'b00000000000000000000000;
mem[130]=23'b00000000000000000000000;
mem[131]=23'b01000100010010100100010;
mem[132]=23'b00000000000000000000000;
mem[133]=23'b00000000000000000000000;
mem[134]=23'b00000000000000000000000;
mem[135]=23'b00000000000000000000000;
mem[136]=23'b00000000000000000000000;
mem[137]=23'b01000110001000101001000;
mem[138]=23'b00000000000000000000000;
mem[139]=23'b00000000000000000000000;
mem[140]=23'b00000000000000000000000;
mem[141]=23'b00000000000000000000000;
mem[142]=23'b00000000000000000000000;
mem[143]=23'b00000000000000000000000;
mem[144]=23'b00000000000000000000000;
mem[145]=23'b00000000000000000000000;
mem[146]=23'b00000000000000000000000;
mem[147]=23'b01000110001100110100100;
mem[148]=23'b00000000000000000000000;
mem[149]=23'b00000000000000000000000;
mem[150]=23'b00000000000000000000000;
mem[151]=23'b00000000000000000000000;
mem[152]=23'b00000000000000000000000;
mem[153]=23'b00000000000000000000000;
mem[154]=23'b00000000000000000000000;
mem[155]=23'b00000000000000000000000;
mem[156]=23'b00000000000000000000000;
mem[157]=23'b00000000000000000000000;
mem[158]=23'b00000000000000000000000;
mem[159]=23'b00000000000000000000000;
mem[160]=23'b00000000000000000000000;
mem[161]=23'b00000000000000000000000;
mem[162]=23'b00000000000000000000000;
mem[163]=23'b00000000000000000000000;
mem[164]=23'b00000000000000000000000;
mem[165]=23'b00000000000000000000000;
mem[166]=23'b00000000000000000000000;
mem[167]=23'b00000000000000000000000;
mem[168]=23'b01000101001000110001001;
mem[169]=23'b01000110001100101000100;
mem[170]=23'b00000000000000000000000;
mem[171]=23'b00000000000000000000000;
mem[172]=23'b00000000000000000000000;
mem[173]=23'b00000000000000000000000;
mem[174]=23'b00000000000000000000000;
mem[175]=23'b00000000000000000000000;
mem[176]=23'b00000000000000000000000;
mem[177]=23'b00000000000000000000000;
mem[178]=23'b00000000000000000000000;
mem[179]=23'b00000000000000000000000;
mem[180]=23'b00000000000000000000000;
mem[181]=23'b00000000000000000000000;
mem[182]=23'b01000100000100011000101;
mem[183]=23'b00000000000000000000000;
mem[184]=23'b00000000000000000000000;
mem[185]=23'b00000000000000000000000;
mem[186]=23'b00000000000000000000000;
mem[187]=23'b00000000000000000000000;
mem[188]=23'b00000000000000000000000;
mem[189]=23'b00000000000000000000000;
mem[190]=23'b00000000000000000000000;
mem[191]=23'b01000011010100110000000;
mem[192]=23'b00000000000000000000000;
mem[193]=23'b00000000000000000000000;
mem[194]=23'b00000000000000000000000;
mem[195]=23'b00000000000000000000000;
mem[196]=23'b00000000000000000000000;
mem[197]=23'b00000000000000000000000;
mem[198]=23'b00000000000000000000000;
mem[199]=23'b01000010001110100100110;
mem[200]=23'b00000000000000000000000;
mem[201]=23'b00000000000000000000000;
mem[202]=23'b00000000000000000000000;
mem[203]=23'b01000100001100110100101;
mem[204]=23'b00000000000000000000000;
mem[205]=23'b00000000000000000000000;
mem[206]=23'b00000000000000000000000;
mem[207]=23'b01000011000110011001100;
mem[208]=23'b00000000000000000000000;
mem[209]=23'b01000111001000101001000;
mem[210]=23'b00000000000000000000000;
mem[211]=23'b01000100000110011001100;
mem[212]=23'b01000100000110011000101;
mem[213]=23'b00000000000000000000000;
mem[214]=23'b01000111001000101001000;
mem[215]=23'b00000000000000000000000;
mem[216]=23'b00000000000000000000000;
mem[217]=23'b00000000000000000000000;
mem[218]=23'b00000000000000000000000;
mem[219]=23'b00000000000000000000000;
mem[220]=23'b00000000000000000000000;
mem[221]=23'b00000000000000000000000;
mem[222]=23'b00000000000000000000000;
mem[223]=23'b00000000000000000000000;
mem[224]=23'b01000010010000110101010;
mem[225]=23'b01000010000110100101101;
mem[226]=23'b00000000000000000000000;
mem[227]=23'b00000000000000000000000;
mem[228]=23'b00000000000000000000000;
mem[229]=23'b00000000000000000000000;
mem[230]=23'b00000000000000000000000;
mem[231]=23'b00000000000000000000000;
mem[232]=23'b00000000000000000000000;
mem[233]=23'b00000000000000000000000;
mem[234]=23'b00000000000000000000000;
mem[235]=23'b00000000000000000000000;
mem[236]=23'b00000000000000000000000;
mem[237]=23'b00000000000000000000000;
mem[238]=23'b00000000000000000000000;
mem[239]=23'b01000011001100101000100;
mem[240]=23'b00000000000000000000000;
mem[241]=23'b00000000000000000000000;
mem[242]=23'b00000000000000000000000;
mem[243]=23'b00000000000000000000000;
mem[244]=23'b00000000000000000000000;
mem[245]=23'b00000000000000000000000;
mem[246]=23'b00000000000000000000000;
mem[247]=23'b00000000000000000000000;
mem[248]=23'b01000010001010100100101;
mem[249]=23'b00000000000000000000000;
mem[250]=23'b00000000000000000000000;
mem[251]=23'b00000000000000000000000;
mem[252]=23'b00000000000000000000000;
mem[253]=23'b01000010000101001001010;
mem[254]=23'b00000000000000000000000;
mem[255]=23'b00000000000000000000000;
mem[256]=23'b00000000000000000000000;
mem[257]=23'b00000000000000000000000;
mem[258]=23'b00000000000000000000000;
mem[259]=23'b00000000000000000000000;
mem[260]=23'b00000000000000000000000;
mem[261]=23'b00000000000000000000000;
mem[262]=23'b00000000000000000000000;
mem[263]=23'b00000000000000000000000;
mem[264]=23'b00000000000000000000000;
mem[265]=23'b00000000000000000000000;
mem[266]=23'b00000000000000000000000;
mem[267]=23'b00000000000000000000000;
mem[268]=23'b00000000000000000000000;
mem[269]=23'b00000000000000000000000;
mem[270]=23'b00000000000000000000000;
mem[271]=23'b00000000000000000000000;
mem[272]=23'b00000000000000000000000;
mem[273]=23'b00000000000000000000000;
mem[274]=23'b00000000000000000000000;
mem[275]=23'b00000000000000000000000;
mem[276]=23'b00000000000000000000000;
mem[277]=23'b00000000000000000000000;
mem[278]=23'b00000000000000000000000;
mem[279]=23'b00000000000000000000000;
mem[280]=23'b01000001000110100101101;
mem[281]=23'b00000000000000000000000;
mem[282]=23'b01000010010100111100000;
mem[283]=23'b00000000000000000000000;
mem[284]=23'b00000000000000000000000;
mem[285]=23'b01000001000110100100100;
mem[286]=23'b01000001010100001100000;
mem[287]=23'b00000000000000000000000;
mem[288]=23'b01000011000111000000111;
mem[289]=23'b00000000000000000000000;
mem[290]=23'b00000000000000000000000;
mem[291]=23'b00000000000000000000000;
mem[292]=23'b01000110001110101000100;
mem[293]=23'b00000000000000000000000;
mem[294]=23'b00000000000000000000000;
mem[295]=23'b00000000000000000000000;
mem[296]=23'b00000000000000000000000;
mem[297]=23'b01000101000100011000101;
mem[298]=23'b00000000000000000000000;
mem[299]=23'b00000000000000000000000;
mem[300]=23'b00000000000000000000000;
mem[301]=23'b00000000000000000000000;
mem[302]=23'b00000000000000000000000;
mem[303]=23'b01000110001100101101010;
mem[304]=23'b00000000000000000000000;
mem[305]=23'b00000000000000000000000;
mem[306]=23'b01000001001110001100011;
mem[307]=23'b00000000000000000000000;
mem[308]=23'b00000000000000000000000;
mem[309]=23'b00000000000000000000000;
mem[310]=23'b00000000000000000000000;
mem[311]=23'b00000000000000000000000;
mem[312]=23'b00000000000000000000000;
mem[313]=23'b00000000000000000000000;
mem[314]=23'b00000000000000000000000;
mem[315]=23'b00000000000000000000000;
mem[316]=23'b00000000000000000000000;
mem[317]=23'b00000000000000000000000;
mem[318]=23'b00000000000000000000000;
mem[319]=23'b00000000000000000000000;
mem[320]=23'b00000000000000000000000;
mem[321]=23'b00000000000000000000000;
mem[322]=23'b01000011010100010100000;
mem[323]=23'b01000101000110011100110;
mem[324]=23'b00000000000000000000000;
mem[325]=23'b00000000000000000000000;
mem[326]=23'b00000000000000000000000;
mem[327]=23'b00000000000000000000000;
mem[328]=23'b00000000000000000000000;
mem[329]=23'b01000011000101000000110;
mem[330]=23'b01000110001000011000110;
mem[331]=23'b00000000000000000000000;
mem[332]=23'b00000000000000000000000;
mem[333]=23'b00000000000000000000000;
mem[334]=23'b00000000000000000000000;
mem[335]=23'b00000000000000000000000;
mem[336]=23'b00000000000000000000000;
mem[337]=23'b00000000000000000000000;
mem[338]=23'b00000000000000000000000;
mem[339]=23'b00000000000000000000000;
mem[340]=23'b00000000000000000000000;
mem[341]=23'b00000000000000000000000;
mem[342]=23'b00000000000000000000000;
mem[343]=23'b00000000000000000000000;
mem[344]=23'b00000000000000000000000;
mem[345]=23'b00000000000000000000000;
mem[346]=23'b00000000000000000000000;
mem[347]=23'b00000000000000000000000;
mem[348]=23'b00000000000000000000000;
mem[349]=23'b00000000000000000000000;
mem[350]=23'b00000000000000000000000;
mem[351]=23'b00000000000000000000000;
mem[352]=23'b00000000000000000000000;
mem[353]=23'b00000000000000000000000;
mem[354]=23'b00000000000000000000000;
mem[355]=23'b00000000000000000000000;
mem[356]=23'b00000000000000000000000;
mem[357]=23'b00000000000000000000000;
mem[358]=23'b00000000000000000000000;
mem[359]=23'b00000000000000000000000;
mem[360]=23'b00000000000000000000000;
mem[361]=23'b00000000000000000000000;
mem[362]=23'b00000000000000000000000;
mem[363]=23'b00000000000000000000000;
mem[364]=23'b00000000000000000000000;
mem[365]=23'b01000010001111000101010;
mem[366]=23'b01000010010000010000010;
mem[367]=23'b00000000000000000000000;
mem[368]=23'b00000000000000000000000;
mem[369]=23'b00000000000000000000000;
mem[370]=23'b01000010000110100101101;
mem[371]=23'b00000000000000000000000;
mem[372]=23'b01000010000110100101101;
mem[373]=23'b01000010000110100100100;
mem[374]=23'b00000000000000000000000;
mem[375]=23'b00000000000000000000000;
mem[376]=23'b00000000000000000000000;
mem[377]=23'b00000000000000000000000;
mem[378]=23'b00000000000000000000000;
mem[379]=23'b01000010000010010000110;
mem[380]=23'b00000000000000000000000;
mem[381]=23'b00000000000000000000000;
mem[382]=23'b00000000000000000000000;
mem[383]=23'b00000000000000000000000;
mem[384]=23'b00000000000000000000000;
mem[385]=23'b01000101000110101001001;
mem[386]=23'b01000110001000101101001;
mem[387]=23'b00000000000000000000000;
mem[388]=23'b00000000000000000000000;
mem[389]=23'b00000000000000000000000;
mem[390]=23'b00000000000000000000000;
mem[391]=23'b00000000000000000000000;
mem[392]=23'b00000000000000000000000;
mem[393]=23'b00000000000000000000000;
mem[394]=23'b00000000000000000000000;
mem[395]=23'b00000000000000000000000;
mem[396]=23'b00000000000000000000000;
mem[397]=23'b00000000000000000000000;
mem[398]=23'b00000000000000000000000;
mem[399]=23'b00000000000000000000000;
mem[400]=23'b00000000000000000000000;
mem[401]=23'b01000011000111000000111;
mem[402]=23'b00000000000000000000000;
mem[403]=23'b00000000000000000000000;
mem[404]=23'b00000000000000000000000;
mem[405]=23'b00000000000000000000000;
mem[406]=23'b00000000000000000000000;
mem[407]=23'b00000000000000000000000;
mem[408]=23'b00000000000000000000000;
mem[409]=23'b00000000000000000000000;
mem[410]=23'b00000000000000000000000;
mem[411]=23'b00000000000000000000000;
mem[412]=23'b00000000000000000000000;
mem[413]=23'b00000000000000000000000;
mem[414]=23'b00000000000000000000000;
mem[415]=23'b00000000000000000000000;
mem[416]=23'b00000000000000000000000;
mem[417]=23'b00000000000000000000000;
mem[418]=23'b00000000000000000000000;
mem[419]=23'b01000010010010001100010;
mem[420]=23'b00000000000000000000000;
mem[421]=23'b01000011001010010100101;
mem[422]=23'b00000000000000000000000;
mem[423]=23'b00000000000000000000000;
mem[424]=23'b00000000000000000000000;
mem[425]=23'b00000000000000000000000;
mem[426]=23'b00000000000000000000000;
mem[427]=23'b00000000000000000000000;
mem[428]=23'b00000000000000000000000;
mem[429]=23'b00000000000000000000000;
mem[430]=23'b00000000000000000000000;
mem[431]=23'b00000000000000000000000;
mem[432]=23'b00000000000000000000000;
mem[433]=23'b00000000000000000000000;
mem[434]=23'b00000000000000000000000;
mem[435]=23'b00000000000000000000000;
mem[436]=23'b00000000000000000000000;
mem[437]=23'b00000000000000000000000;
mem[438]=23'b00000000000000000000000;
mem[439]=23'b00000000000000000000000;
mem[440]=23'b00000000000000000000000;
mem[441]=23'b00000000000000000000000;
mem[442]=23'b01000011000101000100101;
mem[443]=23'b00000000000000000000000;
mem[444]=23'b00000000000000000000000;
mem[445]=23'b00000000000000000000000;
mem[446]=23'b00000000000000000000000;
mem[447]=23'b00000000000000000000000;
mem[448]=23'b00000000000000000000000;
mem[449]=23'b00000000000000000000000;
mem[450]=23'b00000000000000000000000;
mem[451]=23'b00000000000000000000000;
mem[452]=23'b00000000000000000000000;
mem[453]=23'b00000000000000000000000;
mem[454]=23'b00000000000000000000000;
mem[455]=23'b00000000000000000000000;
mem[456]=23'b01000001000010011100111;
mem[457]=23'b01000010010010110100010;
mem[458]=23'b01000001000010011100111;
mem[459]=23'b00000000000000000000000;
mem[460]=23'b00000000000000000000000;
mem[461]=23'b00000000000000000000000;
mem[462]=23'b00000000000000000000000;
mem[463]=23'b00000000000000000000000;
mem[464]=23'b00000000000000000000000;
mem[465]=23'b01000010000110100101001;
mem[466]=23'b00000000000000000000000;
mem[467]=23'b01000010000101000101011;
mem[468]=23'b00000000000000000000000;
mem[469]=23'b00000000000000000000000;
mem[470]=23'b01000010000101000100111;
mem[471]=23'b00000000000000000000000;
mem[472]=23'b00000000000000000000000;
mem[473]=23'b00000000000000000000000;
mem[474]=23'b00000000000000000000000;
mem[475]=23'b00000000000000000000000;
mem[476]=23'b00000000000000000000000;
mem[477]=23'b00000000000000000000000;
mem[478]=23'b00000000000000000000000;
mem[479]=23'b00000000000000000000000;
mem[480]=23'b00000000000000000000000;
mem[481]=23'b00000000000000000000000;
mem[482]=23'b00000000000000000000000;
mem[483]=23'b00000000000000000000000;
mem[484]=23'b00000000000000000000000;
mem[485]=23'b00000000000000000000000;
mem[486]=23'b00000000000000000000000;
mem[487]=23'b00000000000000000000000;
mem[488]=23'b00000000000000000000000;
mem[489]=23'b00000000000000000000000;
mem[490]=23'b00000000000000000000000;
mem[491]=23'b00000000000000000000000;
mem[492]=23'b00000000000000000000000;
mem[493]=23'b00000000000000000000000;
mem[494]=23'b00000000000000000000000;
mem[495]=23'b01000010001111000000011;
mem[496]=23'b01000001000111000001001;
mem[497]=23'b00000000000000000000000;
mem[498]=23'b00000000000000000000000;
mem[499]=23'b00000000000000000000000;
mem[500]=23'b00000000000000000000000;
mem[501]=23'b00000000000000000000000;
mem[502]=23'b00000000000000000000000;
mem[503]=23'b00000000000000000000000;
mem[504]=23'b00000000000000000000000;
mem[505]=23'b00000000000000000000000;
mem[506]=23'b00000000000000000000000;
mem[507]=23'b00000000000000000000000;
mem[508]=23'b00000000000000000000000;
mem[509]=23'b00000000000000000000000;
mem[510]=23'b01000100001110101001010;
mem[511]=23'b00000000000000000000000;
mem[512]=23'b01000110001100101001001;
mem[513]=23'b00000000000000000000000;
mem[514]=23'b00000000000000000000000;
mem[515]=23'b00000000000000000000000;
mem[516]=23'b00000000000000000000000;
mem[517]=23'b00000000000000000000000;
mem[518]=23'b00000000000000000000000;
mem[519]=23'b00000000000000000000000;
mem[520]=23'b01000001000110011101000;
mem[521]=23'b00000000000000000000000;
mem[522]=23'b00000000000000000000000;
mem[523]=23'b00000000000000000000000;
mem[524]=23'b01000010010000110101001;
mem[525]=23'b00000000000000000000000;
mem[526]=23'b00000000000000000000000;
mem[527]=23'b00000000000000000000000;
mem[528]=23'b00000000000000000000000;
mem[529]=23'b00000000000000000000000;
mem[530]=23'b00000000000000000000000;
mem[531]=23'b00000000000000000000000;
mem[532]=23'b00000000000000000000000;
mem[533]=23'b00000000000000000000000;
mem[534]=23'b00000000000000000000000;
mem[535]=23'b00000000000000000000000;
mem[536]=23'b00000000000000000000000;
mem[537]=23'b00000000000000000000000;
mem[538]=23'b00000000000000000000000;
mem[539]=23'b00000000000000000000000;
mem[540]=23'b00000000000000000000000;
mem[541]=23'b00000000000000000000000;
mem[542]=23'b00000000000000000000000;
mem[543]=23'b00000000000000000000000;
mem[544]=23'b00000000000000000000000;
mem[545]=23'b00000000000000000000000;
mem[546]=23'b00000000000000000000000;
mem[547]=23'b00000000000000000000000;
mem[548]=23'b00000000000000000000000;
mem[549]=23'b00000000000000000000000;
mem[550]=23'b01000111010000101001010;
mem[551]=23'b01001001000100101110000;
mem[552]=23'b00000000000000000000000;
mem[553]=23'b01001001000100101110000;
mem[554]=23'b00000000000000000000000;
mem[555]=23'b00000000000000000000000;
mem[556]=23'b00000000000000000000000;
mem[557]=23'b00000000000000000000000;
mem[558]=23'b00000000000000000000000;
mem[559]=23'b00000000000000000000000;
mem[560]=23'b00000000000000000000000;
mem[561]=23'b00000000000000000000000;
mem[562]=23'b00000000000000000000000;
mem[563]=23'b00000000000000000000000;
mem[564]=23'b00000000000000000000000;
mem[565]=23'b01000100001010100100101;
mem[566]=23'b01000010001100100101010;
mem[567]=23'b00000000000000000000000;
mem[568]=23'b01000010000110100101001;
mem[569]=23'b00000000000000000000000;
mem[570]=23'b01000010000111001001001;
mem[571]=23'b00000000000000000000000;
mem[572]=23'b00000000000000000000000;
mem[573]=23'b00000000000000000000000;
mem[574]=23'b00000000000000000000000;
mem[575]=23'b00000000000000000000000;
mem[576]=23'b00000000000000000000000;
mem[577]=23'b00000000000000000000000;
mem[578]=23'b00000000000000000000000;
mem[579]=23'b00000000000000000000000;
mem[580]=23'b00000000000000000000000;
mem[581]=23'b00000000000000000000000;
mem[582]=23'b00000000000000000000000;
mem[583]=23'b00000000000000000000000;
mem[584]=23'b00000000000000000000000;
mem[585]=23'b00000000000000000000000;
mem[586]=23'b00000000000000000000000;
mem[587]=23'b00000000000000000000000;
mem[588]=23'b00000000000000000000000;
mem[589]=23'b00000000000000000000000;
mem[590]=23'b00000000000000000000000;
mem[591]=23'b00000000000000000000000;
mem[592]=23'b00000000000000000000000;
mem[593]=23'b00000000000000000000000;
mem[594]=23'b00000000000000000000000;
mem[595]=23'b00000000000000000000000;
mem[596]=23'b00000000000000000000000;
mem[597]=23'b00000000000000000000000;
mem[598]=23'b00000000000000000000000;
mem[599]=23'b00000000000000000000000;
mem[600]=23'b01000001000010101101011;
mem[601]=23'b00000000000000000000000;
mem[602]=23'b00000000000000000000000;
mem[603]=23'b00000000000000000000000;
mem[604]=23'b00000000000000000000000;
mem[605]=23'b00000000000000000000000;
mem[606]=23'b01000001000010101101011;
mem[607]=23'b00000000000000000000000;
mem[608]=23'b00000000000000000000000;
mem[609]=23'b00000000000000000000000;
mem[610]=23'b00000000000000000000000;
mem[611]=23'b00000000000000000000000;
mem[612]=23'b00000000000000000000000;
mem[613]=23'b00000000000000000000000;
mem[614]=23'b00000000000000000000000;
mem[615]=23'b01000101000110011000011;
mem[616]=23'b00000000000000000000000;
mem[617]=23'b00000000000000000000000;
mem[618]=23'b00000000000000000000000;
mem[619]=23'b00000000000000000000000;
mem[620]=23'b00000000000000000000000;
mem[621]=23'b00000000000000000000000;
mem[622]=23'b01000001000010101101011;
mem[623]=23'b01000001000010101101000;
mem[624]=23'b00000000000000000000000;
mem[625]=23'b00000000000000000000000;
mem[626]=23'b00000000000000000000000;
mem[627]=23'b00000000000000000000000;
mem[628]=23'b01000101001010110000101;
mem[629]=23'b01000001001001001100111;
mem[630]=23'b00000000000000000000000;
mem[631]=23'b00000000000000000000000;
mem[632]=23'b00000000000000000000000;
mem[633]=23'b00000000000000000000000;
mem[634]=23'b00000000000000000000000;
mem[635]=23'b01000001000011000001000;
mem[636]=23'b00000000000000000000000;
mem[637]=23'b00000000000000000000000;
mem[638]=23'b00000000000000000000000;
mem[639]=23'b00000000000000000000000;
mem[640]=23'b00000000000000000000000;
mem[641]=23'b00000000000000000000000;
mem[642]=23'b00000000000000000000000;
mem[643]=23'b00000000000000000000000;
mem[644]=23'b00000000000000000000000;
mem[645]=23'b00000000000000000000000;
mem[646]=23'b00000000000000000000000;
mem[647]=23'b00000000000000000000000;
mem[648]=23'b00000000000000000000000;
mem[649]=23'b00000000000000000000000;
mem[650]=23'b00000000000000000000000;
mem[651]=23'b01000101000010110001001;
mem[652]=23'b00000000000000000000000;
mem[653]=23'b00000000000000000000000;
mem[654]=23'b00000000000000000000000;
mem[655]=23'b00000000000000000000000;
mem[656]=23'b00000000000000000000000;
mem[657]=23'b00000000000000000000000;
mem[658]=23'b00000000000000000000000;
mem[659]=23'b00000000000000000000000;
mem[660]=23'b00000000000000000000000;
mem[661]=23'b00000000000000000000000;
mem[662]=23'b00000000000000000000000;
mem[663]=23'b00000000000000000000000;
mem[664]=23'b00000000000000000000000;
mem[665]=23'b00000000000000000000000;
mem[666]=23'b01001001000010101010010;
mem[667]=23'b00000000000000000000000;
mem[668]=23'b01001001000010101010010;
mem[669]=23'b01000011000101000100011;
mem[670]=23'b00000000000000000000000;
mem[671]=23'b01000101000110111100011;
mem[672]=23'b00000000000000000000000;
mem[673]=23'b00000000000000000000000;
mem[674]=23'b00000000000000000000000;
mem[675]=23'b01000011010010101001010;
mem[676]=23'b00000000000000000000000;
mem[677]=23'b00000000000000000000000;
mem[678]=23'b00000000000000000000000;
mem[679]=23'b00000000000000000000000;
mem[680]=23'b00000000000000000000000;
mem[681]=23'b00000000000000000000000;
mem[682]=23'b00000000000000000000000;
mem[683]=23'b01000010000100100101101;
mem[684]=23'b01000010000100100100101;
mem[685]=23'b00000000000000000000000;
mem[686]=23'b00000000000000000000000;
mem[687]=23'b01000110001010101100110;
mem[688]=23'b00000000000000000000000;
mem[689]=23'b00000000000000000000000;
mem[690]=23'b00000000000000000000000;
mem[691]=23'b00000000000000000000000;
mem[692]=23'b00000000000000000000000;
mem[693]=23'b00000000000000000000000;
mem[694]=23'b00000000000000000000000;
mem[695]=23'b00000000000000000000000;
mem[696]=23'b00000000000000000000000;
mem[697]=23'b00000000000000000000000;
mem[698]=23'b00000000000000000000000;
mem[699]=23'b00000000000000000000000;
mem[700]=23'b00000000000000000000000;
mem[701]=23'b00000000000000000000000;
mem[702]=23'b00000000000000000000000;
mem[703]=23'b00000000000000000000000;
mem[704]=23'b00000000000000000000000;
mem[705]=23'b00000000000000000000000;
mem[706]=23'b00000000000000000000000;
mem[707]=23'b00000000000000000000000;
mem[708]=23'b00000000000000000000000;
mem[709]=23'b01000110001000110000111;
mem[710]=23'b01000110001000110001001;
mem[711]=23'b00000000000000000000000;
mem[712]=23'b00000000000000000000000;
mem[713]=23'b00000000000000000000000;
mem[714]=23'b00000000000000000000000;
mem[715]=23'b00000000000000000000000;
mem[716]=23'b00000000000000000000000;
mem[717]=23'b00000000000000000000000;
mem[718]=23'b00000000000000000000000;
mem[719]=23'b00000000000000000000000;
mem[720]=23'b00000000000000000000000;
mem[721]=23'b00000000000000000000000;
mem[722]=23'b00000000000000000000000;
mem[723]=23'b01000011000101000001000;
mem[724]=23'b00000000000000000000000;
mem[725]=23'b00000000000000000000000;
mem[726]=23'b01000001010100001101010;
mem[727]=23'b00000000000000000000000;
mem[728]=23'b00000000000000000000000;
mem[729]=23'b00000000000000000000000;
mem[730]=23'b00000000000000000000000;
mem[731]=23'b01000100000111000001110;
mem[732]=23'b01000011001011000001001;
mem[733]=23'b00000000000000000000000;
mem[734]=23'b00000000000000000000000;
mem[735]=23'b00000000000000000000000;
mem[736]=23'b00000000000000000000000;
mem[737]=23'b00000000000000000000000;
mem[738]=23'b00000000000000000000000;
mem[739]=23'b00000000000000000000000;
mem[740]=23'b00000000000000000000000;
mem[741]=23'b00000000000000000000000;
mem[742]=23'b00000000000000000000000;
mem[743]=23'b00000000000000000000000;
mem[744]=23'b00000000000000000000000;
mem[745]=23'b00000000000000000000000;
mem[746]=23'b00000000000000000000000;
mem[747]=23'b00000000000000000000000;
mem[748]=23'b01000011000111000100011;
mem[749]=23'b00000000000000000000000;
mem[750]=23'b00000000000000000000000;
mem[751]=23'b00000000000000000000000;
mem[752]=23'b00000000000000000000000;
mem[753]=23'b00000000000000000000000;
mem[754]=23'b00000000000000000000000;
mem[755]=23'b00000000000000000000000;
mem[756]=23'b00000000000000000000000;
mem[757]=23'b00000000000000000000000;
mem[758]=23'b00000000000000000000000;
mem[759]=23'b00000000000000000000000;
mem[760]=23'b01000110001100101001001;
mem[761]=23'b00000000000000000000000;
mem[762]=23'b00000000000000000000000;
mem[763]=23'b00000000000000000000000;
mem[764]=23'b00000000000000000000000;
mem[765]=23'b00000000000000000000000;
mem[766]=23'b00000000000000000000000;
mem[767]=23'b00000000000000000000000;
mem[768]=23'b00000000000000000000000;
mem[769]=23'b01000011010010110100001;
mem[770]=23'b00000000000000000000000;
mem[771]=23'b00000000000000000000000;
mem[772]=23'b00000000000000000000000;
mem[773]=23'b00000000000000000000000;
mem[774]=23'b01000110001100011100111;
mem[775]=23'b01000010000010011001010;
mem[776]=23'b01000001001010101000101;
mem[777]=23'b00000000000000000000000;
mem[778]=23'b00000000000000000000000;
mem[779]=23'b00000000000000000000000;
mem[780]=23'b00000000000000000000000;
mem[781]=23'b01000010000110100101001;
mem[782]=23'b00000000000000000000000;
mem[783]=23'b00000000000000000000000;
mem[784]=23'b00000000000000000000000;
mem[785]=23'b00000000000000000000000;
mem[786]=23'b00000000000000000000000;
mem[787]=23'b00000000000000000000000;
mem[788]=23'b00000000000000000000000;
mem[789]=23'b00000000000000000000000;
mem[790]=23'b00000000000000000000000;
mem[791]=23'b00000000000000000000000;
mem[792]=23'b00000000000000000000000;
mem[793]=23'b00000000000000000000000;
mem[794]=23'b01000011000101000100110;
mem[795]=23'b00000000000000000000000;
mem[796]=23'b00000000000000000000000;
mem[797]=23'b01000100000110010001110;
mem[798]=23'b00000000000000000000000;
mem[799]=23'b00000000000000000000000;
mem[800]=23'b01000110001000011001010;
mem[801]=23'b01000101000010010101110;
mem[802]=23'b01000011001000011001001;
mem[803]=23'b01000101000110010101110;
mem[804]=23'b00000000000000000000000;
mem[805]=23'b00000000000000000000000;
mem[806]=23'b00000000000000000000000;
mem[807]=23'b01000010001110111100011;
mem[808]=23'b00000000000000000000000;
mem[809]=23'b00000000000000000000000;
mem[810]=23'b00000000000000000000000;
mem[811]=23'b00000000000000000000000;
mem[812]=23'b00000000000000000000000;
mem[813]=23'b01000101001100100100100;
mem[814]=23'b00000000000000000000000;
mem[815]=23'b01000100000101000001000;
mem[816]=23'b00000000000000000000000;
mem[817]=23'b00000000000000000000000;
mem[818]=23'b00000000000000000000000;
mem[819]=23'b00000000000000000000000;
mem[820]=23'b00000000000000000000000;
mem[821]=23'b00000000000000000000000;
mem[822]=23'b00000000000000000000000;
mem[823]=23'b00000000000000000000000;
mem[824]=23'b00000000000000000000000;
mem[825]=23'b00000000000000000000000;
mem[826]=23'b00000000000000000000000;
mem[827]=23'b01000100000110010101110;
mem[828]=23'b01000100000110010100011;
mem[829]=23'b01000011010010010100001;
mem[830]=23'b00000000000000000000000;
mem[831]=23'b01000011000100010101101;
mem[832]=23'b00000000000000000000000;
mem[833]=23'b00000000000000000000000;
mem[834]=23'b00000000000000000000000;
mem[835]=23'b01000011000100010101101;
mem[836]=23'b01000011000100010100101;
mem[837]=23'b00000000000000000000000;
mem[838]=23'b00000000000000000000000;
mem[839]=23'b00000000000000000000000;
mem[840]=23'b00000000000000000000000;
mem[841]=23'b00000000000000000000000;
mem[842]=23'b01000010000101001001000;
mem[843]=23'b00000000000000000000000;
mem[844]=23'b00000000000000000000000;
mem[845]=23'b00000000000000000000000;
mem[846]=23'b00000000000000000000000;
mem[847]=23'b00000000000000000000000;
mem[848]=23'b00000000000000000000000;
mem[849]=23'b00000000000000000000000;
mem[850]=23'b00000000000000000000000;
mem[851]=23'b00000000000000000000000;
mem[852]=23'b00000000000000000000000;
mem[853]=23'b00000000000000000000000;
mem[854]=23'b00000000000000000000000;
mem[855]=23'b00000000000000000000000;
mem[856]=23'b00000000000000000000000;
mem[857]=23'b00000000000000000000000;
mem[858]=23'b01000001000010110001000;
mem[859]=23'b00000000000000000000000;
mem[860]=23'b00000000000000000000000;
mem[861]=23'b00000000000000000000000;
mem[862]=23'b00000000000000000000000;
mem[863]=23'b00000000000000000000000;
mem[864]=23'b00000000000000000000000;
mem[865]=23'b00000000000000000000000;
mem[866]=23'b00000000000000000000000;
mem[867]=23'b00000000000000000000000;
mem[868]=23'b00000000000000000000000;
mem[869]=23'b00000000000000000000000;
mem[870]=23'b00000000000000000000000;
mem[871]=23'b00000000000000000000000;
mem[872]=23'b00000000000000000000000;
mem[873]=23'b00000000000000000000000;
mem[874]=23'b00000000000000000000000;
mem[875]=23'b01000101000100111101110;
mem[876]=23'b00000000000000000000000;
mem[877]=23'b00000000000000000000000;
mem[878]=23'b01000101000100111100100;
mem[879]=23'b01000011010101000000000;
mem[880]=23'b00000000000000000000000;
mem[881]=23'b01000010010010100100001;
mem[882]=23'b00000000000000000000000;
mem[883]=23'b01000011010000100100010;
mem[884]=23'b00000000000000000000000;
mem[885]=23'b00000000000000000000000;
mem[886]=23'b01000001001000001101001;
mem[887]=23'b00000000000000000000000;
mem[888]=23'b00000000000000000000000;
mem[889]=23'b00000000000000000000000;
mem[890]=23'b00000000000000000000000;
mem[891]=23'b00000000000000000000000;
mem[892]=23'b00000000000000000000000;
mem[893]=23'b00000000000000000000000;
mem[894]=23'b00000000000000000000000;
mem[895]=23'b00000000000000000000000;
mem[896]=23'b00000000000000000000000;
mem[897]=23'b00000000000000000000000;
mem[898]=23'b00000000000000000000000;
mem[899]=23'b00000000000000000000000;
mem[900]=23'b00000000000000000000000;
mem[901]=23'b00000000000000000000000;
mem[902]=23'b00000000000000000000000;
mem[903]=23'b00000000000000000000000;
mem[904]=23'b00000000000000000000000;
mem[905]=23'b00000000000000000000000;
mem[906]=23'b00000000000000000000000;
mem[907]=23'b00000000000000000000000;
mem[908]=23'b00000000000000000000000;
mem[909]=23'b00000000000000000000000;
mem[910]=23'b00000000000000000000000;
mem[911]=23'b00000000000000000000000;
mem[912]=23'b00000000000000000000000;
mem[913]=23'b00000000000000000000000;
mem[914]=23'b00000000000000000000000;
mem[915]=23'b00000000000000000000000;
mem[916]=23'b00000000000000000000000;
mem[917]=23'b01000010000111001001000;
mem[918]=23'b00000000000000000000000;
mem[919]=23'b00000000000000000000000;
mem[920]=23'b01000101001000101100111;
mem[921]=23'b01000101001000101101001;
mem[922]=23'b00000000000000000000000;
mem[923]=23'b00000000000000000000000;
mem[924]=23'b00000000000000000000000;
mem[925]=23'b01000101000010010100101;
mem[926]=23'b00000000000000000000000;
mem[927]=23'b00000000000000000000000;
mem[928]=23'b00000000000000000000000;
mem[929]=23'b00000000000000000000000;
mem[930]=23'b00000000000000000000000;
mem[931]=23'b00000000000000000000000;
mem[932]=23'b00000000000000000000000;
mem[933]=23'b00000000000000000000000;
mem[934]=23'b00000000000000000000000;
mem[935]=23'b00000000000000000000000;
mem[936]=23'b00000000000000000000000;
mem[937]=23'b00000000000000000000000;
mem[938]=23'b00000000000000000000000;
mem[939]=23'b00000000000000000000000;
mem[940]=23'b00000000000000000000000;
mem[941]=23'b00000000000000000000000;
mem[942]=23'b01000011000010010101011;
mem[943]=23'b00000000000000000000000;
mem[944]=23'b00000000000000000000000;
mem[945]=23'b00000000000000000000000;
mem[946]=23'b00000000000000000000000;
mem[947]=23'b00000000000000000000000;
mem[948]=23'b00000000000000000000000;
mem[949]=23'b00000000000000000000000;
mem[950]=23'b00000000000000000000000;
mem[951]=23'b00000000000000000000000;
mem[952]=23'b01000001000100111101011;
mem[953]=23'b00000000000000000000000;
mem[954]=23'b00000000000000000000000;
mem[955]=23'b00000000000000000000000;
mem[956]=23'b00000000000000000000000;
mem[957]=23'b00000000000000000000000;
mem[958]=23'b00000000000000000000000;
mem[959]=23'b00000000000000000000000;
mem[960]=23'b00000000000000000000000;
mem[961]=23'b00000000000000000000000;
mem[962]=23'b00000000000000000000000;
mem[963]=23'b00000000000000000000000;
mem[964]=23'b00000000000000000000000;
mem[965]=23'b00000000000000000000000;
mem[966]=23'b00000000000000000000000;
mem[967]=23'b00000000000000000000000;
mem[968]=23'b00000000000000000000000;
mem[969]=23'b00000000000000000000000;
mem[970]=23'b00000000000000000000000;
mem[971]=23'b00000000000000000000000;
mem[972]=23'b00000000000000000000000;
mem[973]=23'b00000000000000000000000;
mem[974]=23'b01000101001100010100101;
mem[975]=23'b00000000000000000000000;
mem[976]=23'b00000000000000000000000;
mem[977]=23'b01000101000010011000100;
mem[978]=23'b00000000000000000000000;
mem[979]=23'b00000000000000000000000;
mem[980]=23'b00000000000000000000000;
mem[981]=23'b00000000000000000000000;
mem[982]=23'b01000010010010111000010;
mem[983]=23'b01000001000010100000110;
mem[984]=23'b00000000000000000000000;
mem[985]=23'b01001001000010101100001;
mem[986]=23'b01000010010010010000001;
mem[987]=23'b00000000000000000000000;
mem[988]=23'b01000010010010111000010;
mem[989]=23'b01000010010010111001001;
mem[990]=23'b00000000000000000000000;
mem[991]=23'b00000000000000000000000;
mem[992]=23'b00000000000000000000000;
mem[993]=23'b00000000000000000000000;
mem[994]=23'b00000000000000000000000;
mem[995]=23'b00000000000000000000000;
mem[996]=23'b01000100000010010001011;
mem[997]=23'b01000110000110111000011;
mem[998]=23'b00000000000000000000000;
mem[999]=23'b00000000000000000000000;
mem[1000]=23'b00000000000000000000000;
mem[1001]=23'b00000000000000000000000;
mem[1002]=23'b00000000000000000000000;
mem[1003]=23'b01000100000100010101010;
mem[1004]=23'b00000000000000000000000;
mem[1005]=23'b00000000000000000000000;
mem[1006]=23'b00000000000000000000000;
mem[1007]=23'b00000000000000000000000;
mem[1008]=23'b00000000000000000000000;
mem[1009]=23'b00000000000000000000000;
mem[1010]=23'b00000000000000000000000;
mem[1011]=23'b00000000000000000000000;
mem[1012]=23'b01000101010010100100001;
mem[1013]=23'b00000000000000000000000;
mem[1014]=23'b00000000000000000000000;
mem[1015]=23'b00000000000000000000000;
mem[1016]=23'b00000000000000000000000;
mem[1017]=23'b00000000000000000000000;
mem[1018]=23'b00000000000000000000000;
mem[1019]=23'b00000000000000000000000;
mem[1020]=23'b00000000000000000000000;
mem[1021]=23'b00000000000000000000000;
mem[1022]=23'b01000100000010011110010;
mem[1023]=23'b01000100000010011100001;
mem[1024]=23'b01000101001110110000011;
mem[1025]=23'b00000000000000000000000;
mem[1026]=23'b00000000000000000000000;
mem[1027]=23'b00000000000000000000000;
mem[1028]=23'b00000000000000000000000;
mem[1029]=23'b00000000000000000000000;
mem[1030]=23'b00000000000000000000000;
mem[1031]=23'b00000000000000000000000;
mem[1032]=23'b00000000000000000000000;
mem[1033]=23'b00000000000000000000000;
mem[1034]=23'b00000000000000000000000;
mem[1035]=23'b01000101000110010100011;
mem[1036]=23'b00000000000000000000000;
mem[1037]=23'b00000000000000000000000;
mem[1038]=23'b00000000000000000000000;
mem[1039]=23'b00000000000000000000000;
mem[1040]=23'b01000001001110110000110;
mem[1041]=23'b01000001000010011001001;
mem[1042]=23'b00000000000000000000000;
mem[1043]=23'b00000000000000000000000;
mem[1044]=23'b00000000000000000000000;
mem[1045]=23'b00000000000000000000000;
mem[1046]=23'b00000000000000000000000;
mem[1047]=23'b00000000000000000000000;
mem[1048]=23'b01000011000101000001000;
mem[1049]=23'b00000000000000000000000;
mem[1050]=23'b00000000000000000000000;
mem[1051]=23'b01000011000010010000110;
mem[1052]=23'b00000000000000000000000;
mem[1053]=23'b00000000000000000000000;
mem[1054]=23'b00000000000000000000000;
mem[1055]=23'b00000000000000000000000;
mem[1056]=23'b01000101001110100101000;
mem[1057]=23'b01000111000110110101011;
mem[1058]=23'b01000111000110110100110;
mem[1059]=23'b00000000000000000000000;
mem[1060]=23'b00000000000000000000000;
mem[1061]=23'b01000010001110010100110;
mem[1062]=23'b00000000000000000000000;
mem[1063]=23'b00000000000000000000000;
mem[1064]=23'b00000000000000000000000;
mem[1065]=23'b00000000000000000000000;
mem[1066]=23'b01000010000110100101000;
mem[1067]=23'b00000000000000000000000;
mem[1068]=23'b00000000000000000000000;
mem[1069]=23'b00000000000000000000000;
mem[1070]=23'b00000000000000000000000;
mem[1071]=23'b00000000000000000000000;
mem[1072]=23'b00000000000000000000000;
mem[1073]=23'b00000000000000000000000;
mem[1074]=23'b00000000000000000000000;
mem[1075]=23'b00000000000000000000000;
mem[1076]=23'b00000000000000000000000;
mem[1077]=23'b00000000000000000000000;
mem[1078]=23'b00000000000000000000000;
mem[1079]=23'b00000000000000000000000;
mem[1080]=23'b00000000000000000000000;
mem[1081]=23'b00000000000000000000000;
mem[1082]=23'b00000000000000000000000;
mem[1083]=23'b00000000000000000000000;
mem[1084]=23'b00000000000000000000000;
mem[1085]=23'b00000000000000000000000;
mem[1086]=23'b00000000000000000000000;
mem[1087]=23'b01000001000100011101010;
mem[1088]=23'b01000001000100011101000;
mem[1089]=23'b00000000000000000000000;
mem[1090]=23'b00000000000000000000000;
mem[1091]=23'b00000000000000000000000;
mem[1092]=23'b00000000000000000000000;
mem[1093]=23'b01000010010010010100010;
mem[1094]=23'b00000000000000000000000;
mem[1095]=23'b00000000000000000000000;
mem[1096]=23'b00000000000000000000000;
mem[1097]=23'b00000000000000000000000;
mem[1098]=23'b00000000000000000000000;
mem[1099]=23'b00000000000000000000000;
mem[1100]=23'b00000000000000000000000;
mem[1101]=23'b00000000000000000000000;
mem[1102]=23'b00000000000000000000000;
mem[1103]=23'b00000000000000000000000;
mem[1104]=23'b00000000000000000000000;
mem[1105]=23'b00000000000000000000000;
mem[1106]=23'b00000000000000000000000;
mem[1107]=23'b00000000000000000000000;
mem[1108]=23'b01000011001000110101010;
mem[1109]=23'b00000000000000000000000;
mem[1110]=23'b00000000000000000000000;
mem[1111]=23'b00000000000000000000000;
mem[1112]=23'b00000000000000000000000;
mem[1113]=23'b00000000000000000000000;
mem[1114]=23'b00000000000000000000000;
mem[1115]=23'b00000000000000000000000;
mem[1116]=23'b00000000000000000000000;
mem[1117]=23'b00000000000000000000000;
mem[1118]=23'b00000000000000000000000;
mem[1119]=23'b00000000000000000000000;
mem[1120]=23'b00000000000000000000000;
mem[1121]=23'b01000001010011001100001;
mem[1122]=23'b00000000000000000000000;
mem[1123]=23'b00000000000000000000000;
mem[1124]=23'b00000000000000000000000;
mem[1125]=23'b00000000000000000000000;
mem[1126]=23'b00000000000000000000000;
mem[1127]=23'b00000000000000000000000;
mem[1128]=23'b00000000000000000000000;
mem[1129]=23'b00000000000000000000000;
mem[1130]=23'b00000000000000000000000;
mem[1131]=23'b00000000000000000000000;
mem[1132]=23'b00000000000000000000000;
mem[1133]=23'b00000000000000000000000;
mem[1134]=23'b00000000000000000000000;
mem[1135]=23'b00000000000000000000000;
mem[1136]=23'b00000000000000000000000;
mem[1137]=23'b00000000000000000000000;
mem[1138]=23'b00000000000000000000000;
mem[1139]=23'b01000001001000010101100;
mem[1140]=23'b01000001001000010100100;
mem[1141]=23'b00000000000000000000000;
mem[1142]=23'b00000000000000000000000;
mem[1143]=23'b00000000000000000000000;
mem[1144]=23'b00000000000000000000000;
mem[1145]=23'b01000100000100100001100;
mem[1146]=23'b01000001000010100000111;
mem[1147]=23'b00000000000000000000000;
mem[1148]=23'b00000000000000000000000;
mem[1149]=23'b00000000000000000000000;
mem[1150]=23'b00000000000000000000000;
mem[1151]=23'b00000000000000000000000;
mem[1152]=23'b00000000000000000000000;
mem[1153]=23'b00000000000000000000000;
mem[1154]=23'b00000000000000000000000;
mem[1155]=23'b00000000000000000000000;
mem[1156]=23'b00000000000000000000000;
mem[1157]=23'b00000000000000000000000;
mem[1158]=23'b00000000000000000000000;
mem[1159]=23'b01000010010000110000010;
mem[1160]=23'b00000000000000000000000;
mem[1161]=23'b00000000000000000000000;
mem[1162]=23'b00000000000000000000000;
mem[1163]=23'b00000000000000000000000;
mem[1164]=23'b01000110001000011001010;
mem[1165]=23'b01000001000010100001101;
mem[1166]=23'b00000000000000000000000;
mem[1167]=23'b00000000000000000000000;
mem[1168]=23'b00000000000000000000000;
mem[1169]=23'b00000000000000000000000;
mem[1170]=23'b00000000000000000000000;
mem[1171]=23'b00000000000000000000000;
mem[1172]=23'b00000000000000000000000;
mem[1173]=23'b00000000000000000000000;
mem[1174]=23'b00000000000000000000000;
mem[1175]=23'b00000000000000000000000;
mem[1176]=23'b00000000000000000000000;
mem[1177]=23'b01000011010100100100000;
mem[1178]=23'b01000001000010011100100;
mem[1179]=23'b01000001000010011101111;
mem[1180]=23'b01000001000010011100100;
mem[1181]=23'b00000000000000000000000;
mem[1182]=23'b01000101010000101001010;
mem[1183]=23'b00000000000000000000000;
mem[1184]=23'b00000000000000000000000;
mem[1185]=23'b00000000000000000000000;
mem[1186]=23'b00000000000000000000000;
mem[1187]=23'b00000000000000000000000;
mem[1188]=23'b00000000000000000000000;
mem[1189]=23'b00000000000000000000000;
mem[1190]=23'b00000000000000000000000;
mem[1191]=23'b00000000000000000000000;
mem[1192]=23'b00000000000000000000000;
mem[1193]=23'b01000010000110100101101;
mem[1194]=23'b00000000000000000000000;
mem[1195]=23'b00000000000000000000000;
mem[1196]=23'b01000011000110010101000;
mem[1197]=23'b01000010000111001001001;
mem[1198]=23'b00000000000000000000000;
mem[1199]=23'b00000000000000000000000;
mem[1200]=23'b00000000000000000000000;
mem[1201]=23'b00000000000000000000000;
mem[1202]=23'b00000000000000000000000;
mem[1203]=23'b01000011000110111000111;
mem[1204]=23'b00000000000000000000000;
mem[1205]=23'b00000000000000000000000;
mem[1206]=23'b00000000000000000000000;
mem[1207]=23'b00000000000000000000000;
mem[1208]=23'b00000000000000000000000;
mem[1209]=23'b00000000000000000000000;
mem[1210]=23'b00000000000000000000000;
mem[1211]=23'b00000000000000000000000;
mem[1212]=23'b00000000000000000000000;
mem[1213]=23'b00000000000000000000000;
mem[1214]=23'b00000000000000000000000;
mem[1215]=23'b00000000000000000000000;
mem[1216]=23'b00000000000000000000000;
mem[1217]=23'b00000000000000000000000;
mem[1218]=23'b00000000000000000000000;
mem[1219]=23'b00000000000000000000000;
mem[1220]=23'b00000000000000000000000;
mem[1221]=23'b00000000000000000000000;
mem[1222]=23'b00000000000000000000000;
mem[1223]=23'b00000000000000000000000;
mem[1224]=23'b00000000000000000000000;
mem[1225]=23'b00000000000000000000000;
mem[1226]=23'b00000000000000000000000;
mem[1227]=23'b00000000000000000000000;
mem[1228]=23'b00000000000000000000000;
mem[1229]=23'b00000000000000000000000;
mem[1230]=23'b00000000000000000000000;
mem[1231]=23'b00000000000000000000000;
mem[1232]=23'b01000110001000011001010;
mem[1233]=23'b00000000000000000000000;
mem[1234]=23'b00000000000000000000000;
mem[1235]=23'b00000000000000000000000;
mem[1236]=23'b00000000000000000000000;
mem[1237]=23'b01000001000110110101001;
mem[1238]=23'b00000000000000000000000;
mem[1239]=23'b01000001000010011101011;
mem[1240]=23'b00000000000000000000000;
mem[1241]=23'b01000001000010011101011;
mem[1242]=23'b00000000000000000000000;
mem[1243]=23'b00000000000000000000000;
mem[1244]=23'b00000000000000000000000;
mem[1245]=23'b00000000000000000000000;
mem[1246]=23'b00000000000000000000000;
mem[1247]=23'b00000000000000000000000;
mem[1248]=23'b00000000000000000000000;
mem[1249]=23'b00000000000000000000000;
mem[1250]=23'b00000000000000000000000;
mem[1251]=23'b00000000000000000000000;
mem[1252]=23'b00000000000000000000000;
mem[1253]=23'b01000001000011000001100;
mem[1254]=23'b00000000000000000000000;
mem[1255]=23'b00000000000000000000000;
mem[1256]=23'b00000000000000000000000;
mem[1257]=23'b00000000000000000000000;
mem[1258]=23'b00000000000000000000000;
mem[1259]=23'b00000000000000000000000;
mem[1260]=23'b01000110000010011100101;
mem[1261]=23'b01000011000111000101011;
mem[1262]=23'b01000011000111000100110;
mem[1263]=23'b00000000000000000000000;
mem[1264]=23'b00000000000000000000000;
mem[1265]=23'b00000000000000000000000;
mem[1266]=23'b00000000000000000000000;
mem[1267]=23'b00000000000000000000000;
mem[1268]=23'b01000001000011000000111;
mem[1269]=23'b01000011001000111000110;
mem[1270]=23'b01000001000010011101000;
mem[1271]=23'b01000011010000010100010;
mem[1272]=23'b00000000000000000000000;
mem[1273]=23'b00000000000000000000000;
mem[1274]=23'b00000000000000000000000;
mem[1275]=23'b00000000000000000000000;
mem[1276]=23'b00000000000000000000000;
mem[1277]=23'b00000000000000000000000;
mem[1278]=23'b01001001000100101100011;
mem[1279]=23'b00000000000000000000000;
mem[1280]=23'b00000000000000000000000;
mem[1281]=23'b00000000000000000000000;
mem[1282]=23'b00000000000000000000000;
mem[1283]=23'b00000000000000000000000;
mem[1284]=23'b00000000000000000000000;
mem[1285]=23'b00000000000000000000000;
mem[1286]=23'b00000000000000000000000;
mem[1287]=23'b01000011001000101001100;
mem[1288]=23'b01000011001000101000100;
mem[1289]=23'b01000101000010011110010;
mem[1290]=23'b00000000000000000000000;
mem[1291]=23'b00000000000000000000000;
mem[1292]=23'b01000001000011000001000;
mem[1293]=23'b00000000000000000000000;
mem[1294]=23'b00000000000000000000000;
mem[1295]=23'b00000000000000000000000;
mem[1296]=23'b00000000000000000000000;
mem[1297]=23'b00000000000000000000000;
mem[1298]=23'b00000000000000000000000;
mem[1299]=23'b00000000000000000000000;
mem[1300]=23'b00000000000000000000000;
mem[1301]=23'b00000000000000000000000;
mem[1302]=23'b01000001000010111001000;
mem[1303]=23'b01000010001110110100100;
mem[1304]=23'b00000000000000000000000;
mem[1305]=23'b01000001000011001101011;
mem[1306]=23'b01000001000011001101000;
mem[1307]=23'b00000000000000000000000;
mem[1308]=23'b00000000000000000000000;
mem[1309]=23'b01000100000101000001000;
mem[1310]=23'b00000000000000000000000;
mem[1311]=23'b00000000000000000000000;
mem[1312]=23'b00000000000000000000000;
mem[1313]=23'b00000000000000000000000;
mem[1314]=23'b00000000000000000000000;
mem[1315]=23'b00000000000000000000000;
mem[1316]=23'b00000000000000000000000;
mem[1317]=23'b00000000000000000000000;
mem[1318]=23'b00000000000000000000000;
mem[1319]=23'b01000001000010110001011;
mem[1320]=23'b00000000000000000000000;
mem[1321]=23'b01000001000010110001011;
mem[1322]=23'b00000000000000000000000;
mem[1323]=23'b01000001000010110001011;
mem[1324]=23'b00000000000000000000000;
mem[1325]=23'b01000001000010110001011;
mem[1326]=23'b01000001000010110001000;
mem[1327]=23'b00000000000000000000000;
mem[1328]=23'b00000000000000000000000;
mem[1329]=23'b00000000000000000000000;
mem[1330]=23'b00000000000000000000000;
mem[1331]=23'b00000000000000000000000;
mem[1332]=23'b00000000000000000000000;
mem[1333]=23'b00000000000000000000000;
mem[1334]=23'b01000100000011000001010;
mem[1335]=23'b01000001000010100001011;
mem[1336]=23'b00000000000000000000000;
mem[1337]=23'b00000000000000000000000;
mem[1338]=23'b00000000000000000000000;
mem[1339]=23'b00000000000000000000000;
mem[1340]=23'b00000000000000000000000;
mem[1341]=23'b00000000000000000000000;
mem[1342]=23'b00000000000000000000000;
mem[1343]=23'b00000000000000000000000;
mem[1344]=23'b00000000000000000000000;
mem[1345]=23'b00000000000000000000000;
mem[1346]=23'b00000000000000000000000;
mem[1347]=23'b01000001000010110101100;
mem[1348]=23'b01000001000010110100111;
mem[1349]=23'b01000001000100101001000;
mem[1350]=23'b01000001000010011100100;
mem[1351]=23'b00000000000000000000000;
mem[1352]=23'b00000000000000000000000;
mem[1353]=23'b00000000000000000000000;
mem[1354]=23'b00000000000000000000000;
mem[1355]=23'b00000000000000000000000;
mem[1356]=23'b01000010000110100100100;
mem[1357]=23'b00000000000000000000000;
mem[1358]=23'b00000000000000000000000;
mem[1359]=23'b00000000000000000000000;
mem[1360]=23'b00000000000000000000000;
mem[1361]=23'b00000000000000000000000;
mem[1362]=23'b00000000000000000000000;
mem[1363]=23'b00000000000000000000000;
mem[1364]=23'b00000000000000000000000;
mem[1365]=23'b00000000000000000000000;
mem[1366]=23'b00000000000000000000000;
mem[1367]=23'b00000000000000000000000;
mem[1368]=23'b00000000000000000000000;
mem[1369]=23'b00000000000000000000000;
mem[1370]=23'b00000000000000000000000;
mem[1371]=23'b00000000000000000000000;
mem[1372]=23'b00000000000000000000000;
mem[1373]=23'b00000000000000000000000;
mem[1374]=23'b00000000000000000000000;
mem[1375]=23'b00000000000000000000000;
mem[1376]=23'b00000000000000000000000;
mem[1377]=23'b00000000000000000000000;
mem[1378]=23'b00000000000000000000000;
mem[1379]=23'b00000000000000000000000;
mem[1380]=23'b00000000000000000000000;
mem[1381]=23'b00000000000000000000000;
mem[1382]=23'b00000000000000000000000;
mem[1383]=23'b00000000000000000000000;
mem[1384]=23'b00000000000000000000000;
mem[1385]=23'b00000000000000000000000;
mem[1386]=23'b00000000000000000000000;
mem[1387]=23'b01000011000100001101010;
mem[1388]=23'b00000000000000000000000;
mem[1389]=23'b01000001001000000101100;
mem[1390]=23'b00000000000000000000000;
mem[1391]=23'b01000101000010110010001;
mem[1392]=23'b01000101000010110000010;
mem[1393]=23'b00000000000000000000000;
mem[1394]=23'b00000000000000000000000;
mem[1395]=23'b00000000000000000000000;
mem[1396]=23'b01000001001000000100100;
mem[1397]=23'b00000000000000000000000;
mem[1398]=23'b00000000000000000000000;
mem[1399]=23'b00000000000000000000000;
mem[1400]=23'b00000000000000000000000;
mem[1401]=23'b00000000000000000000000;
mem[1402]=23'b00000000000000000000000;
mem[1403]=23'b00000000000000000000000;
mem[1404]=23'b00000000000000000000000;
mem[1405]=23'b00000000000000000000000;
mem[1406]=23'b00000000000000000000000;
mem[1407]=23'b00000000000000000000000;
mem[1408]=23'b00000000000000000000000;
mem[1409]=23'b00000000000000000000000;
mem[1410]=23'b00000000000000000000000;
mem[1411]=23'b00000000000000000000000;
mem[1412]=23'b00000000000000000000000;
mem[1413]=23'b01000011010100010100000;
mem[1414]=23'b00000000000000000000000;
mem[1415]=23'b00000000000000000000000;
mem[1416]=23'b00000000000000000000000;
mem[1417]=23'b00000000000000000000000;
mem[1418]=23'b00000000000000000000000;
mem[1419]=23'b01000101000100111110000;
mem[1420]=23'b00000000000000000000000;
mem[1421]=23'b00000000000000000000000;
mem[1422]=23'b01000101000100111100010;
mem[1423]=23'b00000000000000000000000;
mem[1424]=23'b00000000000000000000000;
mem[1425]=23'b00000000000000000000000;
mem[1426]=23'b00000000000000000000000;
mem[1427]=23'b00000000000000000000000;
mem[1428]=23'b00000000000000000000000;
mem[1429]=23'b00000000000000000000000;
mem[1430]=23'b00000000000000000000000;
mem[1431]=23'b00000000000000000000000;
mem[1432]=23'b00000000000000000000000;
mem[1433]=23'b00000000000000000000000;
mem[1434]=23'b00000000000000000000000;
mem[1435]=23'b00000000000000000000000;
mem[1436]=23'b00000000000000000000000;
mem[1437]=23'b00000000000000000000000;
mem[1438]=23'b00000000000000000000000;
mem[1439]=23'b00000000000000000000000;
mem[1440]=23'b00000000000000000000000;
mem[1441]=23'b00000000000000000000000;
mem[1442]=23'b00000000000000000000000;
mem[1443]=23'b00000000000000000000000;
mem[1444]=23'b00000000000000000000000;
mem[1445]=23'b00000000000000000000000;
mem[1446]=23'b00000000000000000000000;
mem[1447]=23'b00000000000000000000000;
mem[1448]=23'b00000000000000000000000;
mem[1449]=23'b01000011000010001101011;
mem[1450]=23'b01000011000010001101000;
mem[1451]=23'b00000000000000000000000;
mem[1452]=23'b00000000000000000000000;
mem[1453]=23'b00000000000000000000000;
mem[1454]=23'b00000000000000000000000;
mem[1455]=23'b01000100010000010000010;
mem[1456]=23'b00000000000000000000000;
mem[1457]=23'b00000000000000000000000;
mem[1458]=23'b00000000000000000000000;
mem[1459]=23'b00000000000000000000000;
mem[1460]=23'b00000000000000000000000;
mem[1461]=23'b00000000000000000000000;
mem[1462]=23'b01000010010000100101001;
mem[1463]=23'b00000000000000000000000;
mem[1464]=23'b00000000000000000000000;
mem[1465]=23'b01000101001110101000100;
mem[1466]=23'b00000000000000000000000;
mem[1467]=23'b00000000000000000000000;
mem[1468]=23'b00000000000000000000000;
mem[1469]=23'b00000000000000000000000;
mem[1470]=23'b00000000000000000000000;
mem[1471]=23'b00000000000000000000000;
mem[1472]=23'b00000000000000000000000;
mem[1473]=23'b00000000000000000000000;
mem[1474]=23'b00000000000000000000000;
mem[1475]=23'b00000000000000000000000;
mem[1476]=23'b00000000000000000000000;
mem[1477]=23'b00000000000000000000000;
mem[1478]=23'b00000000000000000000000;
mem[1479]=23'b00000000000000000000000;
mem[1480]=23'b00000000000000000000000;
mem[1481]=23'b00000000000000000000000;
mem[1482]=23'b00000000000000000000000;
mem[1483]=23'b00000000000000000000000;
mem[1484]=23'b00000000000000000000000;
mem[1485]=23'b00000000000000000000000;
mem[1486]=23'b00000000000000000000000;
mem[1487]=23'b00000000000000000000000;
mem[1488]=23'b00000000000000000000000;
mem[1489]=23'b00000000000000000000000;
mem[1490]=23'b00000000000000000000000;
mem[1491]=23'b01000001001001001101001;
mem[1492]=23'b00000000000000000000000;
mem[1493]=23'b00000000000000000000000;
mem[1494]=23'b00000000000000000000000;
mem[1495]=23'b00000000000000000000000;
mem[1496]=23'b00000000000000000000000;
mem[1497]=23'b01000100001110010100100;
mem[1498]=23'b01001000000100110000100;
mem[1499]=23'b00000000000000000000000;
mem[1500]=23'b01000110001010101101001;
mem[1501]=23'b00000000000000000000000;
mem[1502]=23'b00000000000000000000000;
mem[1503]=23'b01000101000100011101100;
mem[1504]=23'b00000000000000000000000;
mem[1505]=23'b01000001010010000100010;
mem[1506]=23'b01000001010010000101001;
mem[1507]=23'b01000011000101000001101;
mem[1508]=23'b01000011000101000000101;
mem[1509]=23'b00000000000000000000000;
mem[1510]=23'b01000101001010111001010;
mem[1511]=23'b01000001000100010101011;
mem[1512]=23'b00000000000000000000000;
mem[1513]=23'b01000101000100011101100;
mem[1514]=23'b00000000000000000000000;
mem[1515]=23'b00000000000000000000000;
mem[1516]=23'b00000000000000000000000;
mem[1517]=23'b01000101000100011101100;
mem[1518]=23'b01000101000100011100110;
mem[1519]=23'b01000001000100010101011;
mem[1520]=23'b00000000000000000000000;
mem[1521]=23'b01000001000100010101011;
mem[1522]=23'b00000000000000000000000;
mem[1523]=23'b01000001000100010101011;
mem[1524]=23'b01000001000100010100111;
mem[1525]=23'b01000110000010011001101;
mem[1526]=23'b00000000000000000000000;
mem[1527]=23'b00000000000000000000000;
mem[1528]=23'b00000000000000000000000;
mem[1529]=23'b00000000000000000000000;
mem[1530]=23'b00000000000000000000000;
mem[1531]=23'b01000010000110100101000;
mem[1532]=23'b00000000000000000000000;
mem[1533]=23'b00000000000000000000000;
mem[1534]=23'b00000000000000000000000;
mem[1535]=23'b01000101000100011100110;
mem[1536]=23'b00000000000000000000000;
mem[1537]=23'b00000000000000000000000;
mem[1538]=23'b00000000000000000000000;
mem[1539]=23'b00000000000000000000000;
mem[1540]=23'b00000000000000000000000;
mem[1541]=23'b00000000000000000000000;
mem[1542]=23'b00000000000000000000000;
mem[1543]=23'b00000000000000000000000;
mem[1544]=23'b00000000000000000000000;
mem[1545]=23'b00000000000000000000000;
mem[1546]=23'b00000000000000000000000;
mem[1547]=23'b00000000000000000000000;
mem[1548]=23'b00000000000000000000000;
mem[1549]=23'b01000101001000010100100;
mem[1550]=23'b00000000000000000000000;
mem[1551]=23'b00000000000000000000000;
mem[1552]=23'b00000000000000000000000;
mem[1553]=23'b00000000000000000000000;
mem[1554]=23'b00000000000000000000000;
mem[1555]=23'b00000000000000000000000;
mem[1556]=23'b00000000000000000000000;
mem[1557]=23'b00000000000000000000000;
mem[1558]=23'b00000000000000000000000;
mem[1559]=23'b00000000000000000000000;
mem[1560]=23'b00000000000000000000000;
mem[1561]=23'b00000000000000000000000;
mem[1562]=23'b00000000000000000000000;
mem[1563]=23'b00000000000000000000000;
mem[1564]=23'b00000000000000000000000;
mem[1565]=23'b00000000000000000000000;
mem[1566]=23'b00000000000000000000000;
mem[1567]=23'b00000000000000000000000;
mem[1568]=23'b00000000000000000000000;
mem[1569]=23'b00000000000000000000000;
mem[1570]=23'b00000000000000000000000;
mem[1571]=23'b00000000000000000000000;
mem[1572]=23'b00000000000000000000000;
mem[1573]=23'b00000000000000000000000;
mem[1574]=23'b00000000000000000000000;
mem[1575]=23'b00000000000000000000000;
mem[1576]=23'b00000000000000000000000;
mem[1577]=23'b00000000000000000000000;
mem[1578]=23'b00000000000000000000000;
mem[1579]=23'b00000000000000000000000;
mem[1580]=23'b00000000000000000000000;
mem[1581]=23'b00000000000000000000000;
mem[1582]=23'b00000000000000000000000;
mem[1583]=23'b00000000000000000000000;
mem[1584]=23'b00000000000000000000000;
mem[1585]=23'b00000000000000000000000;
mem[1586]=23'b00000000000000000000000;
mem[1587]=23'b00000000000000000000000;
mem[1588]=23'b00000000000000000000000;
mem[1589]=23'b00000000000000000000000;
mem[1590]=23'b00000000000000000000000;
mem[1591]=23'b01000110001100101101010;
mem[1592]=23'b01000100001000110100110;
mem[1593]=23'b00000000000000000000000;
mem[1594]=23'b00000000000000000000000;
mem[1595]=23'b00000000000000000000000;
mem[1596]=23'b00000000000000000000000;
mem[1597]=23'b00000000000000000000000;
mem[1598]=23'b00000000000000000000000;
mem[1599]=23'b01000010000100111001001;
mem[1600]=23'b01000001000010110001010;
mem[1601]=23'b00000000000000000000000;
mem[1602]=23'b01000001000010110001010;
mem[1603]=23'b00000000000000000000000;
mem[1604]=23'b01000001000010110001010;
mem[1605]=23'b01000001000010110001001;
mem[1606]=23'b00000000000000000000000;
mem[1607]=23'b00000000000000000000000;
mem[1608]=23'b00000000000000000000000;
mem[1609]=23'b00000000000000000000000;
mem[1610]=23'b01000001000100000101010;
mem[1611]=23'b00000000000000000000000;
mem[1612]=23'b01000100000100111101000;
mem[1613]=23'b00000000000000000000000;
mem[1614]=23'b00000000000000000000000;
mem[1615]=23'b01000110000010110000011;
mem[1616]=23'b00000000000000000000000;
mem[1617]=23'b00000000000000000000000;
mem[1618]=23'b00000000000000000000000;
mem[1619]=23'b00000000000000000000000;
mem[1620]=23'b01000001000100001101001;
mem[1621]=23'b00000000000000000000000;
mem[1622]=23'b00000000000000000000000;
mem[1623]=23'b00000000000000000000000;
mem[1624]=23'b00000000000000000000000;
mem[1625]=23'b00000000000000000000000;
mem[1626]=23'b00000000000000000000000;
mem[1627]=23'b00000000000000000000000;
mem[1628]=23'b00000000000000000000000;
mem[1629]=23'b00000000000000000000000;
mem[1630]=23'b00000000000000000000000;
mem[1631]=23'b00000000000000000000000;
mem[1632]=23'b01000001000110001001001;
mem[1633]=23'b00000000000000000000000;
mem[1634]=23'b01000001000100110101000;
mem[1635]=23'b01000001001010101000110;
mem[1636]=23'b00000000000000000000000;
mem[1637]=23'b00000000000000000000000;
mem[1638]=23'b00000000000000000000000;
mem[1639]=23'b00000000000000000000000;
mem[1640]=23'b00000000000000000000000;
mem[1641]=23'b01000001001000100001001;
mem[1642]=23'b00000000000000000000000;
mem[1643]=23'b00000000000000000000000;
mem[1644]=23'b00000000000000000000000;
mem[1645]=23'b00000000000000000000000;
mem[1646]=23'b00000000000000000000000;
mem[1647]=23'b00000000000000000000000;
mem[1648]=23'b00000000000000000000000;
mem[1649]=23'b00000000000000000000000;
mem[1650]=23'b00000000000000000000000;
mem[1651]=23'b00000000000000000000000;
mem[1652]=23'b00000000000000000000000;
mem[1653]=23'b00000000000000000000000;
mem[1654]=23'b01000100000110100101001;
mem[1655]=23'b01000100000110100101000;
mem[1656]=23'b00000000000000000000000;
mem[1657]=23'b00000000000000000000000;
mem[1658]=23'b00000000000000000000000;
mem[1659]=23'b00000000000000000000000;
mem[1660]=23'b00000000000000000000000;
mem[1661]=23'b00000000000000000000000;
mem[1662]=23'b00000000000000000000000;
mem[1663]=23'b00000000000000000000000;
mem[1664]=23'b00000000000000000000000;
mem[1665]=23'b00000000000000000000000;
mem[1666]=23'b00000000000000000000000;
mem[1667]=23'b00000000000000000000000;
mem[1668]=23'b00000000000000000000000;
mem[1669]=23'b00000000000000000000000;
mem[1670]=23'b00000000000000000000000;
mem[1671]=23'b00000000000000000000000;
mem[1672]=23'b01000101000110110101101;
mem[1673]=23'b00000000000000000000000;
mem[1674]=23'b01000001000010110001100;
mem[1675]=23'b00000000000000000000000;
mem[1676]=23'b00000000000000000000000;
mem[1677]=23'b00000000000000000000000;
mem[1678]=23'b00000000000000000000000;
mem[1679]=23'b00000000000000000000000;
mem[1680]=23'b00000000000000000000000;
mem[1681]=23'b01000001000010110000111;
mem[1682]=23'b00000000000000000000000;
mem[1683]=23'b00000000000000000000000;
mem[1684]=23'b01000100000111000001110;
mem[1685]=23'b00000000000000000000000;
mem[1686]=23'b00000000000000000000000;
mem[1687]=23'b00000000000000000000000;
mem[1688]=23'b00000000000000000000000;
mem[1689]=23'b00000000000000000000000;
mem[1690]=23'b01000010001100101100100;
mem[1691]=23'b01000001000111000001000;
mem[1692]=23'b00000000000000000000000;
mem[1693]=23'b01000001010100111001010;
mem[1694]=23'b01000100001100110100100;
mem[1695]=23'b00000000000000000000000;
mem[1696]=23'b00000000000000000000000;
mem[1697]=23'b01000001000010110101010;
mem[1698]=23'b01000010001110110100100;
mem[1699]=23'b00000000000000000000000;
mem[1700]=23'b00000000000000000000000;
mem[1701]=23'b00000000000000000000000;
mem[1702]=23'b01000110000110111001101;
mem[1703]=23'b01000110000110111000100;
mem[1704]=23'b00000000000000000000000;
mem[1705]=23'b01000010001000110101001;
mem[1706]=23'b01000010001001001001010;
mem[1707]=23'b00000000000000000000000;
mem[1708]=23'b00000000000000000000000;
mem[1709]=23'b00000000000000000000000;
mem[1710]=23'b00000000000000000000000;
mem[1711]=23'b00000000000000000000000;
mem[1712]=23'b00000000000000000000000;
mem[1713]=23'b00000000000000000000000;
mem[1714]=23'b00000000000000000000000;
mem[1715]=23'b00000000000000000000000;
mem[1716]=23'b00000000000000000000000;
mem[1717]=23'b00000000000000000000000;
mem[1718]=23'b01000010001011000101000;
mem[1719]=23'b00000000000000000000000;
mem[1720]=23'b00000000000000000000000;
mem[1721]=23'b00000000000000000000000;
mem[1722]=23'b00000000000000000000000;
mem[1723]=23'b00000000000000000000000;
mem[1724]=23'b00000000000000000000000;
mem[1725]=23'b00000000000000000000000;
mem[1726]=23'b00000000000000000000000;
mem[1727]=23'b00000000000000000000000;
mem[1728]=23'b00000000000000000000000;
mem[1729]=23'b00000000000000000000000;
mem[1730]=23'b00000000000000000000000;
mem[1731]=23'b00000000000000000000000;
mem[1732]=23'b00000000000000000000000;
mem[1733]=23'b00000000000000000000000;
mem[1734]=23'b00000000000000000000000;
mem[1735]=23'b00000000000000000000000;
mem[1736]=23'b00000000000000000000000;
mem[1737]=23'b00000000000000000000000;
mem[1738]=23'b00000000000000000000000;
mem[1739]=23'b00000000000000000000000;
mem[1740]=23'b01000011001100010100110;
mem[1741]=23'b00000000000000000000000;
mem[1742]=23'b01000011001110010100100;
mem[1743]=23'b00000000000000000000000;
mem[1744]=23'b00000000000000000000000;
mem[1745]=23'b00000000000000000000000;
mem[1746]=23'b00000000000000000000000;
mem[1747]=23'b00000000000000000000000;
mem[1748]=23'b00000000000000000000000;
mem[1749]=23'b00000000000000000000000;
mem[1750]=23'b00000000000000000000000;
mem[1751]=23'b00000000000000000000000;
mem[1752]=23'b00000000000000000000000;
mem[1753]=23'b00000000000000000000000;
mem[1754]=23'b00000000000000000000000;
mem[1755]=23'b00000000000000000000000;
mem[1756]=23'b00000000000000000000000;
mem[1757]=23'b00000000000000000000000;
mem[1758]=23'b00000000000000000000000;
mem[1759]=23'b00000000000000000000000;
mem[1760]=23'b00000000000000000000000;
mem[1761]=23'b00000000000000000000000;
mem[1762]=23'b00000000000000000000000;
mem[1763]=23'b01000010001100110001010;
mem[1764]=23'b00000000000000000000000;
mem[1765]=23'b00000000000000000000000;
mem[1766]=23'b01000011000100111101001;
mem[1767]=23'b00000000000000000000000;
mem[1768]=23'b00000000000000000000000;
mem[1769]=23'b00000000000000000000000;
mem[1770]=23'b00000000000000000000000;
mem[1771]=23'b00000000000000000000000;
mem[1772]=23'b00000000000000000000000;
mem[1773]=23'b00000000000000000000000;
mem[1774]=23'b00000000000000000000000;
mem[1775]=23'b00000000000000000000000;
mem[1776]=23'b00000000000000000000000;
mem[1777]=23'b00000000000000000000000;
mem[1778]=23'b01000001000010100001100;
mem[1779]=23'b01000001000010100000110;
mem[1780]=23'b00000000000000000000000;
mem[1781]=23'b00000000000000000000000;
mem[1782]=23'b00000000000000000000000;
mem[1783]=23'b00000000000000000000000;
mem[1784]=23'b00000000000000000000000;
mem[1785]=23'b00000000000000000000000;
mem[1786]=23'b00000000000000000000000;
mem[1787]=23'b00000000000000000000000;
mem[1788]=23'b01000110001010100001001;
mem[1789]=23'b00000000000000000000000;
mem[1790]=23'b00000000000000000000000;
mem[1791]=23'b00000000000000000000000;
mem[1792]=23'b00000000000000000000000;
mem[1793]=23'b01000001000100011101000;
mem[1794]=23'b00000000000000000000000;
mem[1795]=23'b00000000000000000000000;
mem[1796]=23'b00000000000000000000000;
mem[1797]=23'b00000000000000000000000;
mem[1798]=23'b00000000000000000000000;
mem[1799]=23'b00000000000000000000000;
mem[1800]=23'b00000000000000000000000;
mem[1801]=23'b01000010001011001000111;
mem[1802]=23'b01000011001010100100101;
mem[1803]=23'b00000000000000000000000;
mem[1804]=23'b00000000000000000000000;
mem[1805]=23'b00000000000000000000000;
mem[1806]=23'b00000000000000000000000;
mem[1807]=23'b00000000000000000000000;
mem[1808]=23'b00000000000000000000000;
mem[1809]=23'b00000000000000000000000;
mem[1810]=23'b00000000000000000000000;
mem[1811]=23'b00000000000000000000000;
mem[1812]=23'b00000000000000000000000;
mem[1813]=23'b00000000000000000000000;
mem[1814]=23'b01000001001000001101000;
mem[1815]=23'b00000000000000000000000;
mem[1816]=23'b00000000000000000000000;
mem[1817]=23'b00000000000000000000000;
mem[1818]=23'b00000000000000000000000;
mem[1819]=23'b00000000000000000000000;
mem[1820]=23'b01000100000011000001110;
mem[1821]=23'b00000000000000000000000;
mem[1822]=23'b01000100000011000001110;
mem[1823]=23'b01000110001000011001010;
mem[1824]=23'b00000000000000000000000;
mem[1825]=23'b00000000000000000000000;
mem[1826]=23'b01000011000111000101101;
mem[1827]=23'b01000001010101001001010;
mem[1828]=23'b01000011000010011001010;
mem[1829]=23'b00000000000000000000000;
mem[1830]=23'b00000000000000000000000;
mem[1831]=23'b00000000000000000000000;
mem[1832]=23'b00000000000000000000000;
mem[1833]=23'b00000000000000000000000;
mem[1834]=23'b00000000000000000000000;
mem[1835]=23'b00000000000000000000000;
mem[1836]=23'b00000000000000000000000;
mem[1837]=23'b00000000000000000000000;
mem[1838]=23'b01000011001101000101000;
mem[1839]=23'b01000010010100111101010;
mem[1840]=23'b01000001001110011000100;
mem[1841]=23'b01000110001010100000110;
mem[1842]=23'b00000000000000000000000;
mem[1843]=23'b00000000000000000000000;
mem[1844]=23'b00000000000000000000000;
mem[1845]=23'b01000001000101000000111;
mem[1846]=23'b00000000000000000000000;
mem[1847]=23'b01000010000101001001010;
mem[1848]=23'b00000000000000000000000;
mem[1849]=23'b00000000000000000000000;
mem[1850]=23'b01000011000111000101101;
mem[1851]=23'b00000000000000000000000;
mem[1852]=23'b01000011000111000101101;
mem[1853]=23'b00000000000000000000000;
mem[1854]=23'b00000000000000000000000;
mem[1855]=23'b01000011000111000100100;
mem[1856]=23'b01000011000101000101000;
mem[1857]=23'b00000000000000000000000;
mem[1858]=23'b00000000000000000000000;
mem[1859]=23'b00000000000000000000000;
mem[1860]=23'b01000011000101000101100;
mem[1861]=23'b01000011000101000100110;
mem[1862]=23'b01000011000011000101101;
mem[1863]=23'b01000011000011000100110;
mem[1864]=23'b00000000000000000000000;
mem[1865]=23'b00000000000000000000000;
mem[1866]=23'b00000000000000000000000;
mem[1867]=23'b00000000000000000000000;
mem[1868]=23'b00000000000000000000000;
mem[1869]=23'b00000000000000000000000;
mem[1870]=23'b01000100000111000001101;
mem[1871]=23'b00000000000000000000000;
mem[1872]=23'b00000000000000000000000;
mem[1873]=23'b00000000000000000000000;
mem[1874]=23'b00000000000000000000000;
mem[1875]=23'b00000000000000000000000;
mem[1876]=23'b00000000000000000000000;
mem[1877]=23'b00000000000000000000000;
mem[1878]=23'b00000000000000000000000;
mem[1879]=23'b00000000000000000000000;
mem[1880]=23'b00000000000000000000000;
mem[1881]=23'b00000000000000000000000;
mem[1882]=23'b01000100000011000001111;
mem[1883]=23'b00000000000000000000000;
mem[1884]=23'b01000001000110111001001;
mem[1885]=23'b00000000000000000000000;
mem[1886]=23'b00000000000000000000000;
mem[1887]=23'b00000000000000000000000;
mem[1888]=23'b00000000000000000000000;
mem[1889]=23'b00000000000000000000000;
mem[1890]=23'b01000100000011000001111;
mem[1891]=23'b01000100000011000000100;
mem[1892]=23'b00000000000000000000000;
mem[1893]=23'b00000000000000000000000;
mem[1894]=23'b01000001001010011000110;
mem[1895]=23'b00000000000000000000000;
mem[1896]=23'b00000000000000000000000;
mem[1897]=23'b01000001000011000100101;
mem[1898]=23'b00000000000000000000000;
mem[1899]=23'b01000001010101001001010;
mem[1900]=23'b00000000000000000000000;
mem[1901]=23'b00000000000000000000000;
mem[1902]=23'b00000000000000000000000;
mem[1903]=23'b01000001000011001100100;
mem[1904]=23'b00000000000000000000000;
mem[1905]=23'b00000000000000000000000;
mem[1906]=23'b00000000000000000000000;
mem[1907]=23'b01000001000110111101010;
mem[1908]=23'b00000000000000000000000;
mem[1909]=23'b00000000000000000000000;
mem[1910]=23'b00000000000000000000000;
mem[1911]=23'b01000010001111000101001;
mem[1912]=23'b01000001001110100000011;
mem[1913]=23'b00000000000000000000000;
mem[1914]=23'b00000000000000000000000;
mem[1915]=23'b00000000000000000000000;
mem[1916]=23'b00000000000000000000000;
mem[1917]=23'b00000000000000000000000;
mem[1918]=23'b00000000000000000000000;
mem[1919]=23'b00000000000000000000000;
mem[1920]=23'b00000000000000000000000;
mem[1921]=23'b00000000000000000000000;
mem[1922]=23'b00000000000000000000000;
mem[1923]=23'b00000000000000000000000;
mem[1924]=23'b00000000000000000000000;
mem[1925]=23'b00000000000000000000000;
mem[1926]=23'b00000000000000000000000;
mem[1927]=23'b00000000000000000000000;
mem[1928]=23'b00000000000000000000000;
mem[1929]=23'b00000000000000000000000;
mem[1930]=23'b00000000000000000000000;
mem[1931]=23'b01001000000010101101110;
mem[1932]=23'b00000000000000000000000;
mem[1933]=23'b00000000000000000000000;
mem[1934]=23'b01000001000101001101000;
mem[1935]=23'b01000101010000100100010;
mem[1936]=23'b00000000000000000000000;
mem[1937]=23'b00000000000000000000000;
mem[1938]=23'b00000000000000000000000;
mem[1939]=23'b00000000000000000000000;
mem[1940]=23'b00000000000000000000000;
mem[1941]=23'b00000000000000000000000;
mem[1942]=23'b00000000000000000000000;
mem[1943]=23'b00000000000000000000000;
mem[1944]=23'b00000000000000000000000;
mem[1945]=23'b00000000000000000000000;
mem[1946]=23'b00000000000000000000000;
mem[1947]=23'b00000000000000000000000;
mem[1948]=23'b00000000000000000000000;
mem[1949]=23'b00000000000000000000000;
mem[1950]=23'b00000000000000000000000;
mem[1951]=23'b00000000000000000000000;
mem[1952]=23'b00000000000000000000000;
mem[1953]=23'b00000000000000000000000;
mem[1954]=23'b00000000000000000000000;
mem[1955]=23'b01000010001010100000101;
mem[1956]=23'b00000000000000000000000;
mem[1957]=23'b01000001000010110101010;
mem[1958]=23'b00000000000000000000000;
mem[1959]=23'b00000000000000000000000;
mem[1960]=23'b00000000000000000000000;
mem[1961]=23'b00000000000000000000000;
mem[1962]=23'b00000000000000000000000;
mem[1963]=23'b00000000000000000000000;
mem[1964]=23'b00000000000000000000000;
mem[1965]=23'b00000000000000000000000;
mem[1966]=23'b00000000000000000000000;
mem[1967]=23'b00000000000000000000000;
mem[1968]=23'b00000000000000000000000;
mem[1969]=23'b01000100001000110100110;
mem[1970]=23'b01000011000100111101001;
mem[1971]=23'b00000000000000000000000;
mem[1972]=23'b01000101000010110001010;
mem[1973]=23'b00000000000000000000000;
mem[1974]=23'b00000000000000000000000;
mem[1975]=23'b00000000000000000000000;
mem[1976]=23'b01000011000111000100100;
mem[1977]=23'b00000000000000000000000;
mem[1978]=23'b00000000000000000000000;
mem[1979]=23'b00000000000000000000000;
mem[1980]=23'b00000000000000000000000;
mem[1981]=23'b00000000000000000000000;
mem[1982]=23'b00000000000000000000000;
mem[1983]=23'b00000000000000000000000;
mem[1984]=23'b00000000000000000000000;
mem[1985]=23'b00000000000000000000000;
mem[1986]=23'b00000000000000000000000;
mem[1987]=23'b01000001000010110101011;
mem[1988]=23'b01000001000010110101000;
mem[1989]=23'b00000000000000000000000;
mem[1990]=23'b00000000000000000000000;
mem[1991]=23'b00000000000000000000000;
mem[1992]=23'b00000000000000000000000;
mem[1993]=23'b00000000000000000000000;
mem[1994]=23'b00000000000000000000000;
mem[1995]=23'b00000000000000000000000;
mem[1996]=23'b00000000000000000000000;
mem[1997]=23'b01000010001101000000100;
mem[1998]=23'b00000000000000000000000;
mem[1999]=23'b00000000000000000000000;
mem[2000]=23'b01000100000100111001010;
mem[2001]=23'b00000000000000000000000;
mem[2002]=23'b00000000000000000000000;
mem[2003]=23'b00000000000000000000000;
mem[2004]=23'b00000000000000000000000;
mem[2005]=23'b00000000000000000000000;
mem[2006]=23'b01000101000010011000011;
mem[2007]=23'b00000000000000000000000;
mem[2008]=23'b00000000000000000000000;
mem[2009]=23'b00000000000000000000000;
mem[2010]=23'b00000000000000000000000;
mem[2011]=23'b01000001000110011001101;
mem[2012]=23'b00000000000000000000000;
mem[2013]=23'b00000000000000000000000;
mem[2014]=23'b00000000000000000000000;
mem[2015]=23'b00000000000000000000000;
mem[2016]=23'b00000000000000000000000;
mem[2017]=23'b00000000000000000000000;
mem[2018]=23'b00000000000000000000000;
mem[2019]=23'b00000000000000000000000;
mem[2020]=23'b00000000000000000000000;
mem[2021]=23'b00000000000000000000000;
mem[2022]=23'b00000000000000000000000;
mem[2023]=23'b00000000000000000000000;
mem[2024]=23'b01000011010000111001010;
mem[2025]=23'b01000001000010100001100;
mem[2026]=23'b00000000000000000000000;
mem[2027]=23'b00000000000000000000000;
mem[2028]=23'b00000000000000000000000;
mem[2029]=23'b00000000000000000000000;
mem[2030]=23'b00000000000000000000000;
mem[2031]=23'b00000000000000000000000;
mem[2032]=23'b00000000000000000000000;
mem[2033]=23'b00000000000000000000000;
mem[2034]=23'b00000000000000000000000;
mem[2035]=23'b01000011000011000101001;
mem[2036]=23'b00000000000000000000000;
mem[2037]=23'b00000000000000000000000;
mem[2038]=23'b00000000000000000000000;
mem[2039]=23'b00000000000000000000000;
mem[2040]=23'b00000000000000000000000;
mem[2041]=23'b00000000000000000000000;
mem[2042]=23'b01000001000010100000110;
mem[2043]=23'b00000000000000000000000;
mem[2044]=23'b00000000000000000000000;
mem[2045]=23'b00000000000000000000000;
mem[2046]=23'b01001000000010101100001;
mem[2047]=23'b00000000000000000000000;
mem[2048]=23'b00000000000000000000000;
mem[2049]=23'b00000000000000000000000;
mem[2050]=23'b00000000000000000000000;
mem[2051]=23'b00000000000000000000000;
mem[2052]=23'b00000000000000000000000;
mem[2053]=23'b00000000000000000000000;
mem[2054]=23'b00000000000000000000000;
mem[2055]=23'b00000000000000000000000;
mem[2056]=23'b01000011010010010001001;
mem[2057]=23'b00000000000000000000000;
mem[2058]=23'b00000000000000000000000;
mem[2059]=23'b00000000000000000000000;
mem[2060]=23'b00000000000000000000000;
mem[2061]=23'b00000000000000000000000;
mem[2062]=23'b00000000000000000000000;
mem[2063]=23'b00000000000000000000000;
mem[2064]=23'b00000000000000000000000;
mem[2065]=23'b00000000000000000000000;
mem[2066]=23'b00000000000000000000000;
mem[2067]=23'b00000000000000000000000;
mem[2068]=23'b00000000000000000000000;
mem[2069]=23'b01000010000110001001101;
mem[2070]=23'b00000000000000000000000;
mem[2071]=23'b00000000000000000000000;
mem[2072]=23'b00000000000000000000000;
mem[2073]=23'b00000000000000000000000;
mem[2074]=23'b00000000000000000000000;
mem[2075]=23'b00000000000000000000000;
mem[2076]=23'b00000000000000000000000;
mem[2077]=23'b00000000000000000000000;
mem[2078]=23'b00000000000000000000000;
mem[2079]=23'b00000000000000000000000;
mem[2080]=23'b00000000000000000000000;
mem[2081]=23'b00000000000000000000000;
mem[2082]=23'b01000001000100011001000;
mem[2083]=23'b00000000000000000000000;
mem[2084]=23'b00000000000000000000000;
mem[2085]=23'b00000000000000000000000;
mem[2086]=23'b00000000000000000000000;
mem[2087]=23'b00000000000000000000000;
mem[2088]=23'b01000010000110001000100;
mem[2089]=23'b00000000000000000000000;
mem[2090]=23'b00000000000000000000000;
mem[2091]=23'b00000000000000000000000;
mem[2092]=23'b00000000000000000000000;
mem[2093]=23'b00000000000000000000000;
mem[2094]=23'b00000000000000000000000;
mem[2095]=23'b01000110000100110001000;
mem[2096]=23'b00000000000000000000000;
mem[2097]=23'b00000000000000000000000;
mem[2098]=23'b00000000000000000000000;
mem[2099]=23'b00000000000000000000000;
mem[2100]=23'b00000000000000000000000;
mem[2101]=23'b00000000000000000000000;
mem[2102]=23'b01000010000101000001001;
mem[2103]=23'b01000011000101000101101;
mem[2104]=23'b00000000000000000000000;
mem[2105]=23'b01000100000010010010000;
mem[2106]=23'b01000100000010010000011;
mem[2107]=23'b00000000000000000000000;
mem[2108]=23'b00000000000000000000000;
mem[2109]=23'b00000000000000000000000;
mem[2110]=23'b00000000000000000000000;
mem[2111]=23'b00000000000000000000000;
mem[2112]=23'b00000000000000000000000;
mem[2113]=23'b00000000000000000000000;
mem[2114]=23'b00000000000000000000000;
mem[2115]=23'b00000000000000000000000;
mem[2116]=23'b00000000000000000000000;
mem[2117]=23'b00000000000000000000000;
mem[2118]=23'b00000000000000000000000;
mem[2119]=23'b00000000000000000000000;
mem[2120]=23'b00000000000000000000000;
mem[2121]=23'b00000000000000000000000;
mem[2122]=23'b00000000000000000000000;
mem[2123]=23'b00000000000000000000000;
mem[2124]=23'b00000000000000000000000;
mem[2125]=23'b00000000000000000000000;
mem[2126]=23'b00000000000000000000000;
mem[2127]=23'b00000000000000000000000;
mem[2128]=23'b00000000000000000000000;
mem[2129]=23'b00000000000000000000000;
mem[2130]=23'b00000000000000000000000;
mem[2131]=23'b00000000000000000000000;
mem[2132]=23'b00000000000000000000000;
mem[2133]=23'b00000000000000000000000;
mem[2134]=23'b01000011001010001100101;
end

always@(posedge clk)
begin
  if (we) begin
    mem[addr] <= din;
  end
end

always @(posedge clk) dout <= mem[addr];

endmodule