library verilog;
use verilog.vl_types.all;
entity UpDown_tb is
end UpDown_tb;
