`timescale 1ns/1ps
module FEAT_RIGHT_ROM(
  addr,
  clk,
  din,
  dout,
  we);

input [11 : 0] addr;
input clk;
input [11 : 0] din;
output reg [11 : 0] dout;
input we;

reg [11:0] mem [0:4095];

initial begin
mem[0]=12'b110101100111;
mem[1]=12'b101111111011;
mem[2]=12'b101000110011;
mem[3]=12'b101101100000;
mem[4]=12'b101010101011;
mem[5]=12'b101001111100;
mem[6]=12'b000101110110;
mem[7]=12'b100110100110;
mem[8]=12'b110010101100;
mem[9]=12'b001101010111;
mem[10]=12'b101000101101;
mem[11]=12'b100101000111;
mem[12]=12'b100101000010;
mem[13]=12'b001000101101;
mem[14]=12'b011110001100;
mem[15]=12'b010010001001;
mem[16]=12'b101101001011;
mem[17]=12'b100110101110;
mem[18]=12'b100100010100;
mem[19]=12'b001001000111;
mem[20]=12'b001000001111;
mem[21]=12'b100111101000;
mem[22]=12'b100100010010;
mem[23]=12'b100101110010;
mem[24]=12'b100100101110;
mem[25]=12'b100101000000;
mem[26]=12'b100100011100;
mem[27]=12'b100110000111;
mem[28]=12'b100011010101;
mem[29]=12'b100011100100;
mem[30]=12'b100111100110;
mem[31]=12'b100011000010;
mem[32]=12'b100100100011;
mem[33]=12'b010101001111;
mem[34]=12'b100011110110;
mem[35]=12'b100111001111;
mem[36]=12'b010110001001;
mem[37]=12'b101100101111;
mem[38]=12'b110001111011;
mem[39]=12'b001000011100;
mem[40]=12'b100111101011;
mem[41]=12'b001100000100;
mem[42]=12'b100101011111;
mem[43]=12'b101000101100;
mem[44]=12'b001101111011;
mem[45]=12'b010011000100;
mem[46]=12'b100101100111;
mem[47]=12'b100001001111;
mem[48]=12'b100101001110;
mem[49]=12'b100100011110;
mem[50]=12'b110000011000;
mem[51]=12'b100011111011;
mem[52]=12'b010000111010;
mem[53]=12'b010001100111;
mem[54]=12'b100100110100;
mem[55]=12'b001110111100;
mem[56]=12'b001101001101;
mem[57]=12'b010011101001;
mem[58]=12'b100111000111;
mem[59]=12'b100110100011;
mem[60]=12'b100010010100;
mem[61]=12'b100011011000;
mem[62]=12'b101101011100;
mem[63]=12'b101000111010;
mem[64]=12'b100010110001;
mem[65]=12'b010100101110;
mem[66]=12'b010010101000;
mem[67]=12'b100001010000;
mem[68]=12'b100011011010;
mem[69]=12'b101100101001;
mem[70]=12'b100011001011;
mem[71]=12'b001111010001;
mem[72]=12'b101100101100;
mem[73]=12'b100010100000;
mem[74]=12'b010011111110;
mem[75]=12'b001011010101;
mem[76]=12'b000111110000;
mem[77]=12'b010101001100;
mem[78]=12'b011100011111;
mem[79]=12'b100110111001;
mem[80]=12'b001000000010;
mem[81]=12'b100100101010;
mem[82]=12'b100100011100;
mem[83]=12'b100101000011;
mem[84]=12'b100011010000;
mem[85]=12'b001011111000;
mem[86]=12'b001110000000;
mem[87]=12'b011001111000;
mem[88]=12'b100010111110;
mem[89]=12'b100011110010;
mem[90]=12'b010000110000;
mem[91]=12'b101001110100;
mem[92]=12'b100011011100;
mem[93]=12'b100011011111;
mem[94]=12'b010011011001;
mem[95]=12'b100100001000;
mem[96]=12'b100010111101;
mem[97]=12'b100010111100;
mem[98]=12'b010001111110;
mem[99]=12'b100011001110;
mem[100]=12'b010101001001;
mem[101]=12'b100010011011;
mem[102]=12'b001110101001;
mem[103]=12'b011011001101;
mem[104]=12'b100010010001;
mem[105]=12'b101111101000;
mem[106]=12'b010000100001;
mem[107]=12'b100010010011;
mem[108]=12'b011101001000;
mem[109]=12'b100010001100;
mem[110]=12'b100011110110;
mem[111]=12'b010001101110;
mem[112]=12'b100111011001;
mem[113]=12'b001011101110;
mem[114]=12'b100100101000;
mem[115]=12'b001111001101;
mem[116]=12'b100101011111;
mem[117]=12'b100101000101;
mem[118]=12'b001111111001;
mem[119]=12'b100011000110;
mem[120]=12'b100110101110;
mem[121]=12'b100010110100;
mem[122]=12'b001111010011;
mem[123]=12'b100110001011;
mem[124]=12'b001010000101;
mem[125]=12'b101011001100;
mem[126]=12'b100011000001;
mem[127]=12'b100001011101;
mem[128]=12'b100111000110;
mem[129]=12'b100010100101;
mem[130]=12'b001110010010;
mem[131]=12'b001111101101;
mem[132]=12'b100010011010;
mem[133]=12'b010100001100;
mem[134]=12'b101010001110;
mem[135]=12'b100011001110;
mem[136]=12'b001100000110;
mem[137]=12'b010101011001;
mem[138]=12'b001111010101;
mem[139]=12'b011001101111;
mem[140]=12'b011101000100;
mem[141]=12'b100010010010;
mem[142]=12'b101101111101;
mem[143]=12'b010001110111;
mem[144]=12'b011001100010;
mem[145]=12'b100001111011;
mem[146]=12'b100001011110;
mem[147]=12'b100010111001;
mem[148]=12'b011100011010;
mem[149]=12'b100011001000;
mem[150]=12'b011011001101;
mem[151]=12'b001110101011;
mem[152]=12'b011001101111;
mem[153]=12'b001001110101;
mem[154]=12'b100001100010;
mem[155]=12'b011011101011;
mem[156]=12'b001001011001;
mem[157]=12'b100101101111;
mem[158]=12'b001011010001;
mem[159]=12'b100011110100;
mem[160]=12'b100100101011;
mem[161]=12'b100011111111;
mem[162]=12'b100100001001;
mem[163]=12'b100011001110;
mem[164]=12'b100100110111;
mem[165]=12'b010111011011;
mem[166]=12'b100101111000;
mem[167]=12'b100111100100;
mem[168]=12'b010100000100;
mem[169]=12'b001100010001;
mem[170]=12'b101010100001;
mem[171]=12'b100100100010;
mem[172]=12'b100011111001;
mem[173]=12'b011101010100;
mem[174]=12'b010010111001;
mem[175]=12'b110000110000;
mem[176]=12'b001011010110;
mem[177]=12'b100010001011;
mem[178]=12'b100110100100;
mem[179]=12'b100010000100;
mem[180]=12'b100010000011;
mem[181]=12'b100001010110;
mem[182]=12'b010110010000;
mem[183]=12'b001110011100;
mem[184]=12'b100001010010;
mem[185]=12'b011000011100;
mem[186]=12'b101010011111;
mem[187]=12'b100010011100;
mem[188]=12'b011010111110;
mem[189]=12'b100010011110;
mem[190]=12'b101011111000;
mem[191]=12'b010110001100;
mem[192]=12'b011011100101;
mem[193]=12'b100001011100;
mem[194]=12'b100011000101;
mem[195]=12'b110100010111;
mem[196]=12'b100001100010;
mem[197]=12'b101111001110;
mem[198]=12'b011100100111;
mem[199]=12'b100011011100;
mem[200]=12'b100010000001;
mem[201]=12'b100000111000;
mem[202]=12'b010101100010;
mem[203]=12'b100001000010;
mem[204]=12'b011100101111;
mem[205]=12'b100110010011;
mem[206]=12'b101010100001;
mem[207]=12'b010000000111;
mem[208]=12'b001111010110;
mem[209]=12'b010000001011;
mem[210]=12'b100011100011;
mem[211]=12'b011110011110;
mem[212]=12'b010010001011;
mem[213]=12'b100110011100;
mem[214]=12'b010001010100;
mem[215]=12'b010100111000;
mem[216]=12'b011010111000;
mem[217]=12'b100010110010;
mem[218]=12'b001110110101;
mem[219]=12'b010001010101;
mem[220]=12'b100101101100;
mem[221]=12'b100010101100;
mem[222]=12'b010001011100;
mem[223]=12'b100110100000;
mem[224]=12'b001001001100;
mem[225]=12'b100101111100;
mem[226]=12'b010011010101;
mem[227]=12'b100011011001;
mem[228]=12'b010101100000;
mem[229]=12'b100001011110;
mem[230]=12'b000110100101;
mem[231]=12'b100011100100;
mem[232]=12'b001100000000;
mem[233]=12'b011101111100;
mem[234]=12'b011011101111;
mem[235]=12'b100100001010;
mem[236]=12'b100001100110;
mem[237]=12'b100010110110;
mem[238]=12'b101000000001;
mem[239]=12'b100100011110;
mem[240]=12'b101001101111;
mem[241]=12'b100010101111;
mem[242]=12'b011001011101;
mem[243]=12'b100001011001;
mem[244]=12'b100011001110;
mem[245]=12'b100111001011;
mem[246]=12'b100001010000;
mem[247]=12'b011111010100;
mem[248]=12'b100011000001;
mem[249]=12'b100110110111;
mem[250]=12'b011101100110;
mem[251]=12'b100001111101;
mem[252]=12'b010000100010;
mem[253]=12'b100100101101;
mem[254]=12'b011100110001;
mem[255]=12'b011010011111;
mem[256]=12'b011011101100;
mem[257]=12'b001111111000;
mem[258]=12'b001110110111;
mem[259]=12'b100101001101;
mem[260]=12'b100101100010;
mem[261]=12'b100101000100;
mem[262]=12'b100100000100;
mem[263]=12'b100110110000;
mem[264]=12'b010001011110;
mem[265]=12'b010111010010;
mem[266]=12'b100010110001;
mem[267]=12'b101101001111;
mem[268]=12'b100001111000;
mem[269]=12'b001111111111;
mem[270]=12'b100100100001;
mem[271]=12'b101111010100;
mem[272]=12'b001111110111;
mem[273]=12'b100010001010;
mem[274]=12'b100010000100;
mem[275]=12'b100011011010;
mem[276]=12'b101001111110;
mem[277]=12'b011000011000;
mem[278]=12'b100100100010;
mem[279]=12'b100001101010;
mem[280]=12'b100100101001;
mem[281]=12'b010011011111;
mem[282]=12'b100011101010;
mem[283]=12'b101001101110;
mem[284]=12'b100011110101;
mem[285]=12'b100011100110;
mem[286]=12'b100010001001;
mem[287]=12'b011011000001;
mem[288]=12'b001101110111;
mem[289]=12'b011011110111;
mem[290]=12'b010110100011;
mem[291]=12'b100010001010;
mem[292]=12'b010111101100;
mem[293]=12'b011101010101;
mem[294]=12'b011001100101;
mem[295]=12'b011000001011;
mem[296]=12'b100001001001;
mem[297]=12'b010111101011;
mem[298]=12'b100100010110;
mem[299]=12'b011100101011;
mem[300]=12'b100010000000;
mem[301]=12'b011010011011;
mem[302]=12'b100011111101;
mem[303]=12'b010001011010;
mem[304]=12'b101010110101;
mem[305]=12'b001010011110;
mem[306]=12'b010010110011;
mem[307]=12'b011101000000;
mem[308]=12'b010110111110;
mem[309]=12'b100010110100;
mem[310]=12'b011001110000;
mem[311]=12'b011100010011;
mem[312]=12'b001011100000;
mem[313]=12'b010000110011;
mem[314]=12'b100100101111;
mem[315]=12'b100100000000;
mem[316]=12'b001100100001;
mem[317]=12'b100110010110;
mem[318]=12'b100110111010;
mem[319]=12'b100011101100;
mem[320]=12'b100011010010;
mem[321]=12'b011100101001;
mem[322]=12'b010001000101;
mem[323]=12'b010011001000;
mem[324]=12'b100000101100;
mem[325]=12'b010011111110;
mem[326]=12'b100100010110;
mem[327]=12'b100010001101;
mem[328]=12'b100010100000;
mem[329]=12'b100100011011;
mem[330]=12'b100011000110;
mem[331]=12'b100100110101;
mem[332]=12'b011110010000;
mem[333]=12'b010010110001;
mem[334]=12'b011011010110;
mem[335]=12'b100001010100;
mem[336]=12'b001010101110;
mem[337]=12'b010001110001;
mem[338]=12'b011110110011;
mem[339]=12'b101000101000;
mem[340]=12'b100010010011;
mem[341]=12'b101111011011;
mem[342]=12'b100010101010;
mem[343]=12'b001000011001;
mem[344]=12'b010000100101;
mem[345]=12'b001010001000;
mem[346]=12'b011100001001;
mem[347]=12'b010111101110;
mem[348]=12'b100011100011;
mem[349]=12'b010101110101;
mem[350]=12'b011011110100;
mem[351]=12'b100001001111;
mem[352]=12'b011110011110;
mem[353]=12'b010101110101;
mem[354]=12'b100011100011;
mem[355]=12'b011110000100;
mem[356]=12'b011001011101;
mem[357]=12'b011000100111;
mem[358]=12'b100001111011;
mem[359]=12'b100101010011;
mem[360]=12'b100001101101;
mem[361]=12'b000110100011;
mem[362]=12'b011011111001;
mem[363]=12'b110000101011;
mem[364]=12'b001011111001;
mem[365]=12'b001110111011;
mem[366]=12'b010100111001;
mem[367]=12'b011101000000;
mem[368]=12'b100010101001;
mem[369]=12'b101101101011;
mem[370]=12'b100011000001;
mem[371]=12'b010100000010;
mem[372]=12'b010101111101;
mem[373]=12'b100010111111;
mem[374]=12'b100010001110;
mem[375]=12'b011100110000;
mem[376]=12'b100001011011;
mem[377]=12'b010011001010;
mem[378]=12'b011100100011;
mem[379]=12'b100010011110;
mem[380]=12'b011110101110;
mem[381]=12'b010100110111;
mem[382]=12'b100100101110;
mem[383]=12'b100001011111;
mem[384]=12'b101011110101;
mem[385]=12'b010000001111;
mem[386]=12'b010001111111;
mem[387]=12'b100011011110;
mem[388]=12'b100010110001;
mem[389]=12'b100111110100;
mem[390]=12'b010011001001;
mem[391]=12'b100010101000;
mem[392]=12'b100010010101;
mem[393]=12'b100100101010;
mem[394]=12'b100001101001;
mem[395]=12'b011000101001;
mem[396]=12'b010111010001;
mem[397]=12'b100010011010;
mem[398]=12'b100011101010;
mem[399]=12'b011101000000;
mem[400]=12'b010010110001;
mem[401]=12'b100010000111;
mem[402]=12'b100000110000;
mem[403]=12'b101100110110;
mem[404]=12'b100000101010;
mem[405]=12'b001000010111;
mem[406]=12'b100010110100;
mem[407]=12'b110001001100;
mem[408]=12'b010100101111;
mem[409]=12'b100001011110;
mem[410]=12'b100011010100;
mem[411]=12'b100111001111;
mem[412]=12'b100001110010;
mem[413]=12'b011111000101;
mem[414]=12'b100001101000;
mem[415]=12'b101000001011;
mem[416]=12'b011101010001;
mem[417]=12'b100011000000;
mem[418]=12'b101011010100;
mem[419]=12'b011000010001;
mem[420]=12'b100101100101;
mem[421]=12'b100011101111;
mem[422]=12'b011101011101;
mem[423]=12'b100101110000;
mem[424]=12'b001011100100;
mem[425]=12'b010111110010;
mem[426]=12'b100000111100;
mem[427]=12'b011110010100;
mem[428]=12'b101000010101;
mem[429]=12'b010111101100;
mem[430]=12'b100000101001;
mem[431]=12'b100001000101;
mem[432]=12'b101000011010;
mem[433]=12'b100010011010;
mem[434]=12'b010111011100;
mem[435]=12'b010110101010;
mem[436]=12'b100100010001;
mem[437]=12'b100001010001;
mem[438]=12'b100000001011;
mem[439]=12'b100111110100;
mem[440]=12'b100000111000;
mem[441]=12'b010111110100;
mem[442]=12'b011101111111;
mem[443]=12'b011011001000;
mem[444]=12'b010110011010;
mem[445]=12'b011110010000;
mem[446]=12'b000100110110;
mem[447]=12'b100011011100;
mem[448]=12'b100010010011;
mem[449]=12'b011101110000;
mem[450]=12'b011011110100;
mem[451]=12'b001110110100;
mem[452]=12'b010011000011;
mem[453]=12'b011111000111;
mem[454]=12'b100001011110;
mem[455]=12'b100001010110;
mem[456]=12'b101010001001;
mem[457]=12'b100001010001;
mem[458]=12'b011101110001;
mem[459]=12'b100101110000;
mem[460]=12'b100010010101;
mem[461]=12'b110101001101;
mem[462]=12'b100010010111;
mem[463]=12'b100110001100;
mem[464]=12'b010011100011;
mem[465]=12'b010100001100;
mem[466]=12'b100100011011;
mem[467]=12'b100101111110;
mem[468]=12'b100011000010;
mem[469]=12'b100100010001;
mem[470]=12'b100101011010;
mem[471]=12'b100011010110;
mem[472]=12'b100010011001;
mem[473]=12'b100011001100;
mem[474]=12'b101000011010;
mem[475]=12'b011001111011;
mem[476]=12'b001110110101;
mem[477]=12'b100001100010;
mem[478]=12'b010111100010;
mem[479]=12'b100011011110;
mem[480]=12'b100001111011;
mem[481]=12'b100101000101;
mem[482]=12'b100001110111;
mem[483]=12'b011110011000;
mem[484]=12'b100011101100;
mem[485]=12'b100001110101;
mem[486]=12'b010110010011;
mem[487]=12'b011101111011;
mem[488]=12'b011101110101;
mem[489]=12'b100010001111;
mem[490]=12'b010101000011;
mem[491]=12'b011110011011;
mem[492]=12'b100010010011;
mem[493]=12'b010110101110;
mem[494]=12'b001000000010;
mem[495]=12'b001010011001;
mem[496]=12'b011101010101;
mem[497]=12'b010110010111;
mem[498]=12'b100001000001;
mem[499]=12'b100100111010;
mem[500]=12'b100010001110;
mem[501]=12'b101000111000;
mem[502]=12'b011010010111;
mem[503]=12'b101101010111;
mem[504]=12'b010010100001;
mem[505]=12'b100001011001;
mem[506]=12'b011111111111;
mem[507]=12'b011001110010;
mem[508]=12'b100101100010;
mem[509]=12'b011111011110;
mem[510]=12'b100010001110;
mem[511]=12'b100111001110;
mem[512]=12'b010101111010;
mem[513]=12'b100101010001;
mem[514]=12'b010010010001;
mem[515]=12'b100110001000;
mem[516]=12'b011110010110;
mem[517]=12'b100010001010;
mem[518]=12'b101011000010;
mem[519]=12'b010010001101;
mem[520]=12'b100100100110;
mem[521]=12'b010001111100;
mem[522]=12'b010101001101;
mem[523]=12'b101000001011;
mem[524]=12'b001100111010;
mem[525]=12'b011111001101;
mem[526]=12'b100101101000;
mem[527]=12'b100001110101;
mem[528]=12'b011101010111;
mem[529]=12'b100011000111;
mem[530]=12'b100001101000;
mem[531]=12'b100010111001;
mem[532]=12'b011100101101;
mem[533]=12'b011001000111;
mem[534]=12'b011101010111;
mem[535]=12'b100010010111;
mem[536]=12'b010111101101;
mem[537]=12'b101001010011;
mem[538]=12'b011010000000;
mem[539]=12'b100001111000;
mem[540]=12'b100000111011;
mem[541]=12'b011111000011;
mem[542]=12'b011010100101;
mem[543]=12'b011101001110;
mem[544]=12'b100001001101;
mem[545]=12'b001110000110;
mem[546]=12'b100000011000;
mem[547]=12'b000111100101;
mem[548]=12'b101011101011;
mem[549]=12'b100001011100;
mem[550]=12'b100000100001;
mem[551]=12'b011110101010;
mem[552]=12'b001010000000;
mem[553]=12'b101110010001;
mem[554]=12'b100000101000;
mem[555]=12'b101011010101;
mem[556]=12'b100000100001;
mem[557]=12'b011110110010;
mem[558]=12'b100001100000;
mem[559]=12'b011111011110;
mem[560]=12'b100110111011;
mem[561]=12'b010101000100;
mem[562]=12'b011101011010;
mem[563]=12'b100100111010;
mem[564]=12'b010000110111;
mem[565]=12'b100001110010;
mem[566]=12'b100011010011;
mem[567]=12'b101000100010;
mem[568]=12'b010110010000;
mem[569]=12'b100011101110;
mem[570]=12'b100101111100;
mem[571]=12'b010101011011;
mem[572]=12'b100011010000;
mem[573]=12'b010111101011;
mem[574]=12'b100010110011;
mem[575]=12'b001011011111;
mem[576]=12'b011100011101;
mem[577]=12'b100010001110;
mem[578]=12'b100010000111;
mem[579]=12'b011101010111;
mem[580]=12'b001110100011;
mem[581]=12'b011000011010;
mem[582]=12'b010000010001;
mem[583]=12'b010101110011;
mem[584]=12'b100010101100;
mem[585]=12'b100100001110;
mem[586]=12'b011001001110;
mem[587]=12'b101101100011;
mem[588]=12'b100010000011;
mem[589]=12'b100000110001;
mem[590]=12'b101001010100;
mem[591]=12'b001111000111;
mem[592]=12'b011100101001;
mem[593]=12'b100000101001;
mem[594]=12'b001001110101;
mem[595]=12'b010111001100;
mem[596]=12'b011111000000;
mem[597]=12'b100101010001;
mem[598]=12'b001001001101;
mem[599]=12'b100001110101;
mem[600]=12'b100111001011;
mem[601]=12'b100000010010;
mem[602]=12'b011110101011;
mem[603]=12'b001111111111;
mem[604]=12'b010111101111;
mem[605]=12'b100000100001;
mem[606]=12'b011110100111;
mem[607]=12'b011100110011;
mem[608]=12'b100010101011;
mem[609]=12'b000111110001;
mem[610]=12'b100010011100;
mem[611]=12'b100100100000;
mem[612]=12'b100011100000;
mem[613]=12'b100000100111;
mem[614]=12'b011011100010;
mem[615]=12'b101100101011;
mem[616]=12'b001110100001;
mem[617]=12'b011101000010;
mem[618]=12'b010001100010;
mem[619]=12'b100000011101;
mem[620]=12'b100111001010;
mem[621]=12'b001100111110;
mem[622]=12'b100010110000;
mem[623]=12'b101011011000;
mem[624]=12'b010101111101;
mem[625]=12'b100000000001;
mem[626]=12'b001010001011;
mem[627]=12'b011101101111;
mem[628]=12'b011001000110;
mem[629]=12'b011101101000;
mem[630]=12'b100001010100;
mem[631]=12'b010011100010;
mem[632]=12'b100001000101;
mem[633]=12'b011011000100;
mem[634]=12'b011010000111;
mem[635]=12'b011101010001;
mem[636]=12'b100001001111;
mem[637]=12'b100000010001;
mem[638]=12'b011110011100;
mem[639]=12'b100000011010;
mem[640]=12'b100100010000;
mem[641]=12'b100011110000;
mem[642]=12'b011110110011;
mem[643]=12'b100001110101;
mem[644]=12'b100101111010;
mem[645]=12'b000100011011;
mem[646]=12'b011111100100;
mem[647]=12'b100101101101;
mem[648]=12'b100010100010;
mem[649]=12'b100000011011;
mem[650]=12'b011011001010;
mem[651]=12'b011101000011;
mem[652]=12'b010011010111;
mem[653]=12'b010000010111;
mem[654]=12'b100101100001;
mem[655]=12'b001001110001;
mem[656]=12'b011111010011;
mem[657]=12'b011100111001;
mem[658]=12'b100010100100;
mem[659]=12'b100000011110;
mem[660]=12'b100010100100;
mem[661]=12'b011101011010;
mem[662]=12'b011100110011;
mem[663]=12'b100001111111;
mem[664]=12'b011110011100;
mem[665]=12'b100010111000;
mem[666]=12'b011110111000;
mem[667]=12'b100001000000;
mem[668]=12'b101101110100;
mem[669]=12'b011101100100;
mem[670]=12'b001111101011;
mem[671]=12'b101000111010;
mem[672]=12'b100011000110;
mem[673]=12'b010001010010;
mem[674]=12'b100010011110;
mem[675]=12'b010111110011;
mem[676]=12'b101100001000;
mem[677]=12'b011001000100;
mem[678]=12'b101101101101;
mem[679]=12'b100110111110;
mem[680]=12'b100110010100;
mem[681]=12'b100100011101;
mem[682]=12'b100011011001;
mem[683]=12'b100100010011;
mem[684]=12'b100010011111;
mem[685]=12'b100011001100;
mem[686]=12'b010001101011;
mem[687]=12'b100001101010;
mem[688]=12'b011010000100;
mem[689]=12'b100010101010;
mem[690]=12'b010110011010;
mem[691]=12'b010101110101;
mem[692]=12'b100010001001;
mem[693]=12'b100011011011;
mem[694]=12'b100001100101;
mem[695]=12'b101010010001;
mem[696]=12'b100001110101;
mem[697]=12'b011110011001;
mem[698]=12'b100000101000;
mem[699]=12'b100101101000;
mem[700]=12'b111010001011;
mem[701]=12'b100011101100;
mem[702]=12'b101010000111;
mem[703]=12'b011001011100;
mem[704]=12'b010111000100;
mem[705]=12'b001011011111;
mem[706]=12'b100000101110;
mem[707]=12'b101010010010;
mem[708]=12'b011100011001;
mem[709]=12'b011001111100;
mem[710]=12'b010100111100;
mem[711]=12'b011111110110;
mem[712]=12'b010110110010;
mem[713]=12'b100101001110;
mem[714]=12'b010110000011;
mem[715]=12'b101111110100;
mem[716]=12'b101000111110;
mem[717]=12'b010110110000;
mem[718]=12'b100100111100;
mem[719]=12'b100001110111;
mem[720]=12'b001010101110;
mem[721]=12'b101101010110;
mem[722]=12'b001101110101;
mem[723]=12'b100001100110;
mem[724]=12'b011010110111;
mem[725]=12'b100010110000;
mem[726]=12'b010000000101;
mem[727]=12'b011111000010;
mem[728]=12'b100010100001;
mem[729]=12'b011101001111;
mem[730]=12'b010001111011;
mem[731]=12'b011101101010;
mem[732]=12'b100001101000;
mem[733]=12'b011010001000;
mem[734]=12'b100101001010;
mem[735]=12'b100001001010;
mem[736]=12'b010110000111;
mem[737]=12'b100110000010;
mem[738]=12'b101100111101;
mem[739]=12'b011000000111;
mem[740]=12'b100010111011;
mem[741]=12'b100000111111;
mem[742]=12'b010001110111;
mem[743]=12'b011110011100;
mem[744]=12'b011010001100;
mem[745]=12'b100001110100;
mem[746]=12'b011101110001;
mem[747]=12'b011100110100;
mem[748]=12'b011101010000;
mem[749]=12'b100001001010;
mem[750]=12'b100001001111;
mem[751]=12'b011111000011;
mem[752]=12'b100011010100;
mem[753]=12'b011010111011;
mem[754]=12'b011101001100;
mem[755]=12'b001110011100;
mem[756]=12'b100001000000;
mem[757]=12'b101010110100;
mem[758]=12'b100001100110;
mem[759]=12'b011111110010;
mem[760]=12'b100000011001;
mem[761]=12'b011011000111;
mem[762]=12'b100011001011;
mem[763]=12'b100100010000;
mem[764]=12'b011100100100;
mem[765]=12'b100001011010;
mem[766]=12'b100000000010;
mem[767]=12'b001000001101;
mem[768]=12'b101111001000;
mem[769]=12'b100011010100;
mem[770]=12'b010111100101;
mem[771]=12'b011110001011;
mem[772]=12'b011000001010;
mem[773]=12'b100001010001;
mem[774]=12'b011000100100;
mem[775]=12'b100100110101;
mem[776]=12'b100001000100;
mem[777]=12'b101001010101;
mem[778]=12'b100110011101;
mem[779]=12'b100011001010;
mem[780]=12'b010111111101;
mem[781]=12'b010110000000;
mem[782]=12'b100101110100;
mem[783]=12'b010010011001;
mem[784]=12'b100010110000;
mem[785]=12'b100100101111;
mem[786]=12'b010110001010;
mem[787]=12'b100010101111;
mem[788]=12'b100010010000;
mem[789]=12'b100100011110;
mem[790]=12'b010101100011;
mem[791]=12'b101000000011;
mem[792]=12'b100000110101;
mem[793]=12'b011010100101;
mem[794]=12'b100101001001;
mem[795]=12'b100001010011;
mem[796]=12'b010110111100;
mem[797]=12'b100110000001;
mem[798]=12'b100000100100;
mem[799]=12'b101011110010;
mem[800]=12'b010111111111;
mem[801]=12'b011000101010;
mem[802]=12'b100010001011;
mem[803]=12'b100110110010;
mem[804]=12'b100110011110;
mem[805]=12'b001011110001;
mem[806]=12'b011100001110;
mem[807]=12'b100011110001;
mem[808]=12'b001101001100;
mem[809]=12'b011010110101;
mem[810]=12'b011001100111;
mem[811]=12'b100010110101;
mem[812]=12'b011001001111;
mem[813]=12'b011010110101;
mem[814]=12'b011101011110;
mem[815]=12'b010010101110;
mem[816]=12'b101110110001;
mem[817]=12'b100010101010;
mem[818]=12'b100011110111;
mem[819]=12'b100001111000;
mem[820]=12'b011101100101;
mem[821]=12'b100010101100;
mem[822]=12'b100000001111;
mem[823]=12'b100011111011;
mem[824]=12'b100101111011;
mem[825]=12'b010111110111;
mem[826]=12'b010011000010;
mem[827]=12'b011110111000;
mem[828]=12'b101001000011;
mem[829]=12'b010101111100;
mem[830]=12'b100000000101;
mem[831]=12'b011110000100;
mem[832]=12'b101001001100;
mem[833]=12'b100110101011;
mem[834]=12'b010100101011;
mem[835]=12'b100001010010;
mem[836]=12'b011000011010;
mem[837]=12'b011110000000;
mem[838]=12'b101000001111;
mem[839]=12'b010101001001;
mem[840]=12'b100000000010;
mem[841]=12'b011011101011;
mem[842]=12'b100010110111;
mem[843]=12'b101011011000;
mem[844]=12'b010111000111;
mem[845]=12'b010100110011;
mem[846]=12'b101010101010;
mem[847]=12'b011000110110;
mem[848]=12'b101110101110;
mem[849]=12'b100010111110;
mem[850]=12'b100000100100;
mem[851]=12'b011111100111;
mem[852]=12'b110010011011;
mem[853]=12'b010001100101;
mem[854]=12'b011001110111;
mem[855]=12'b011110110100;
mem[856]=12'b101100111111;
mem[857]=12'b100001111100;
mem[858]=12'b011110000000;
mem[859]=12'b100011101010;
mem[860]=12'b100001101100;
mem[861]=12'b100010011110;
mem[862]=12'b101111101010;
mem[863]=12'b100011110010;
mem[864]=12'b011101111011;
mem[865]=12'b010101001011;
mem[866]=12'b010101001011;
mem[867]=12'b100110111001;
mem[868]=12'b100101100001;
mem[869]=12'b011010111011;
mem[870]=12'b011001100110;
mem[871]=12'b011011010000;
mem[872]=12'b010101011100;
mem[873]=12'b101101101111;
mem[874]=12'b100000100010;
mem[875]=12'b100000001000;
mem[876]=12'b100011010110;
mem[877]=12'b100010011111;
mem[878]=12'b110000000001;
mem[879]=12'b100011011100;
mem[880]=12'b011100111111;
mem[881]=12'b100011000001;
mem[882]=12'b100101000110;
mem[883]=12'b011100010111;
mem[884]=12'b101000101110;
mem[885]=12'b100101110110;
mem[886]=12'b011000110111;
mem[887]=12'b010111111101;
mem[888]=12'b100011111011;
mem[889]=12'b100001001011;
mem[890]=12'b100100010111;
mem[891]=12'b001111001110;
mem[892]=12'b011100100101;
mem[893]=12'b100001100110;
mem[894]=12'b010101101111;
mem[895]=12'b011111000000;
mem[896]=12'b010110000110;
mem[897]=12'b100001001101;
mem[898]=12'b100100001100;
mem[899]=12'b011111101111;
mem[900]=12'b100000001101;
mem[901]=12'b010001101000;
mem[902]=12'b100001010111;
mem[903]=12'b011100110111;
mem[904]=12'b101110111011;
mem[905]=12'b011010010000;
mem[906]=12'b001000001001;
mem[907]=12'b100001000011;
mem[908]=12'b011101111110;
mem[909]=12'b011110101001;
mem[910]=12'b100001011010;
mem[911]=12'b100001100010;
mem[912]=12'b001111100001;
mem[913]=12'b011110011101;
mem[914]=12'b100001101011;
mem[915]=12'b100111111100;
mem[916]=12'b101100011011;
mem[917]=12'b100101110000;
mem[918]=12'b100001111011;
mem[919]=12'b010011110111;
mem[920]=12'b010110001100;
mem[921]=12'b010101000101;
mem[922]=12'b011000101001;
mem[923]=12'b100111010111;
mem[924]=12'b100010000100;
mem[925]=12'b011000100110;
mem[926]=12'b100100110101;
mem[927]=12'b100011000001;
mem[928]=12'b100111000111;
mem[929]=12'b100001001101;
mem[930]=12'b011110001111;
mem[931]=12'b100001101010;
mem[932]=12'b011001000101;
mem[933]=12'b100111001010;
mem[934]=12'b100010001011;
mem[935]=12'b011100100000;
mem[936]=12'b100010001100;
mem[937]=12'b010101100000;
mem[938]=12'b000101001100;
mem[939]=12'b100001001101;
mem[940]=12'b001110111100;
mem[941]=12'b011011011111;
mem[942]=12'b100011100111;
mem[943]=12'b101010000110;
mem[944]=12'b010111100000;
mem[945]=12'b011101101101;
mem[946]=12'b010001010100;
mem[947]=12'b001111101011;
mem[948]=12'b100011100000;
mem[949]=12'b011010010000;
mem[950]=12'b011111001010;
mem[951]=12'b100001110101;
mem[952]=12'b011101100010;
mem[953]=12'b001011101001;
mem[954]=12'b100001011111;
mem[955]=12'b100111100001;
mem[956]=12'b011011100001;
mem[957]=12'b100000000000;
mem[958]=12'b101011000000;
mem[959]=12'b100001001000;
mem[960]=12'b100111110010;
mem[961]=12'b011100001110;
mem[962]=12'b100010111110;
mem[963]=12'b011111111110;
mem[964]=12'b100001110000;
mem[965]=12'b011101010000;
mem[966]=12'b011010100110;
mem[967]=12'b011011110110;
mem[968]=12'b101011001100;
mem[969]=12'b001100000011;
mem[970]=12'b100001101010;
mem[971]=12'b010001110001;
mem[972]=12'b011110000010;
mem[973]=12'b100001000101;
mem[974]=12'b100001001011;
mem[975]=12'b100010010100;
mem[976]=12'b011011111111;
mem[977]=12'b011010111100;
mem[978]=12'b011110011000;
mem[979]=12'b010101111010;
mem[980]=12'b101000100001;
mem[981]=12'b011011000011;
mem[982]=12'b100010110000;
mem[983]=12'b011110000100;
mem[984]=12'b100010100011;
mem[985]=12'b011110011000;
mem[986]=12'b100011101100;
mem[987]=12'b101100111101;
mem[988]=12'b011000011001;
mem[989]=12'b001010110011;
mem[990]=12'b101000110000;
mem[991]=12'b011100101110;
mem[992]=12'b010011001000;
mem[993]=12'b100000100000;
mem[994]=12'b100001101001;
mem[995]=12'b011100110000;
mem[996]=12'b010001000001;
mem[997]=12'b101101010110;
mem[998]=12'b011000000011;
mem[999]=12'b100001100001;
mem[1000]=12'b100101001001;
mem[1001]=12'b011000110010;
mem[1002]=12'b100100010111;
mem[1003]=12'b011011101000;
mem[1004]=12'b011011110011;
mem[1005]=12'b011101000010;
mem[1006]=12'b011010011110;
mem[1007]=12'b100100100101;
mem[1008]=12'b100001011000;
mem[1009]=12'b011000011100;
mem[1010]=12'b011011001001;
mem[1011]=12'b011010110010;
mem[1012]=12'b100001011100;
mem[1013]=12'b011110001011;
mem[1014]=12'b010101001110;
mem[1015]=12'b011100100010;
mem[1016]=12'b010111010110;
mem[1017]=12'b001010000010;
mem[1018]=12'b101000001111;
mem[1019]=12'b011001001111;
mem[1020]=12'b100000000101;
mem[1021]=12'b100000110100;
mem[1022]=12'b100100110101;
mem[1023]=12'b011101001010;
mem[1024]=12'b001101111111;
mem[1025]=12'b001101011000;
mem[1026]=12'b101101011111;
mem[1027]=12'b100000111111;
mem[1028]=12'b011100011010;
mem[1029]=12'b011101100100;
mem[1030]=12'b100010110111;
mem[1031]=12'b100000110110;
mem[1032]=12'b101001000000;
mem[1033]=12'b100000000110;
mem[1034]=12'b100001000111;
mem[1035]=12'b011101111100;
mem[1036]=12'b000110101001;
mem[1037]=12'b100011011001;
mem[1038]=12'b100001110001;
mem[1039]=12'b011001001010;
mem[1040]=12'b011110011100;
mem[1041]=12'b100011011011;
mem[1042]=12'b100001001111;
mem[1043]=12'b100011110011;
mem[1044]=12'b011110000111;
mem[1045]=12'b011000011000;
mem[1046]=12'b100111001111;
mem[1047]=12'b100010101111;
mem[1048]=12'b011010110100;
mem[1049]=12'b011100100111;
mem[1050]=12'b011110000011;
mem[1051]=12'b011001010000;
mem[1052]=12'b011000110010;
mem[1053]=12'b100110001110;
mem[1054]=12'b010000010011;
mem[1055]=12'b100010011110;
mem[1056]=12'b010110100101;
mem[1057]=12'b100100111001;
mem[1058]=12'b100011011011;
mem[1059]=12'b100011100000;
mem[1060]=12'b011101010011;
mem[1061]=12'b011000111111;
mem[1062]=12'b100001101101;
mem[1063]=12'b010111110001;
mem[1064]=12'b011010010100;
mem[1065]=12'b100010000110;
mem[1066]=12'b011000000101;
mem[1067]=12'b011110000111;
mem[1068]=12'b100011100110;
mem[1069]=12'b100001011000;
mem[1070]=12'b010011100110;
mem[1071]=12'b010010011110;
mem[1072]=12'b100101011101;
mem[1073]=12'b010010010111;
mem[1074]=12'b011101101111;
mem[1075]=12'b100001100101;
mem[1076]=12'b100101111101;
mem[1077]=12'b010100000010;
mem[1078]=12'b100000100010;
mem[1079]=12'b010111111100;
mem[1080]=12'b101111100101;
mem[1081]=12'b100001110010;
mem[1082]=12'b010110010010;
mem[1083]=12'b011111100100;
mem[1084]=12'b001110011010;
mem[1085]=12'b100001101100;
mem[1086]=12'b101101010001;
mem[1087]=12'b100100010001;
mem[1088]=12'b100100100111;
mem[1089]=12'b010011111011;
mem[1090]=12'b100001101110;
mem[1091]=12'b100001100100;
mem[1092]=12'b011110000010;
mem[1093]=12'b100010100111;
mem[1094]=12'b011100010001;
mem[1095]=12'b011001011011;
mem[1096]=12'b100001101100;
mem[1097]=12'b011110011001;
mem[1098]=12'b010101100000;
mem[1099]=12'b000111100000;
mem[1100]=12'b001000111010;
mem[1101]=12'b011111011111;
mem[1102]=12'b100000010100;
mem[1103]=12'b100110101101;
mem[1104]=12'b011101011101;
mem[1105]=12'b100001011100;
mem[1106]=12'b010101100110;
mem[1107]=12'b100001111100;
mem[1108]=12'b011001011011;
mem[1109]=12'b011010000000;
mem[1110]=12'b101100000101;
mem[1111]=12'b010111001100;
mem[1112]=12'b100000000000;
mem[1113]=12'b001100110100;
mem[1114]=12'b101000101111;
mem[1115]=12'b011111001001;
mem[1116]=12'b100010000001;
mem[1117]=12'b100011110111;
mem[1118]=12'b100000110001;
mem[1119]=12'b100001010100;
mem[1120]=12'b011101011111;
mem[1121]=12'b100001100011;
mem[1122]=12'b011000001100;
mem[1123]=12'b011101100001;
mem[1124]=12'b100101011010;
mem[1125]=12'b011010110010;
mem[1126]=12'b100001100000;
mem[1127]=12'b100010010010;
mem[1128]=12'b001111001101;
mem[1129]=12'b100000010100;
mem[1130]=12'b011101111100;
mem[1131]=12'b100010000100;
mem[1132]=12'b100100010110;
mem[1133]=12'b100001111001;
mem[1134]=12'b101111110000;
mem[1135]=12'b011110011010;
mem[1136]=12'b100000000110;
mem[1137]=12'b011111010101;
mem[1138]=12'b100010001101;
mem[1139]=12'b011110101111;
mem[1140]=12'b110000110010;
mem[1141]=12'b011010110100;
mem[1142]=12'b100010100011;
mem[1143]=12'b100010101110;
mem[1144]=12'b011101000111;
mem[1145]=12'b100001001101;
mem[1146]=12'b011110011001;
mem[1147]=12'b100001001000;
mem[1148]=12'b100000111011;
mem[1149]=12'b011101110111;
mem[1150]=12'b100111010001;
mem[1151]=12'b100001001111;
mem[1152]=12'b010011011111;
mem[1153]=12'b101100000101;
mem[1154]=12'b100000000111;
mem[1155]=12'b100001100011;
mem[1156]=12'b011110010011;
mem[1157]=12'b001111010010;
mem[1158]=12'b011100011000;
mem[1159]=12'b011010100011;
mem[1160]=12'b000011111010;
mem[1161]=12'b100010101101;
mem[1162]=12'b100001111011;
mem[1163]=12'b011111101110;
mem[1164]=12'b010010010110;
mem[1165]=12'b101000011011;
mem[1166]=12'b011111111000;
mem[1167]=12'b011110001000;
mem[1168]=12'b011111110111;
mem[1169]=12'b100010011010;
mem[1170]=12'b100011011010;
mem[1171]=12'b011110111000;
mem[1172]=12'b011001110110;
mem[1173]=12'b100001101010;
mem[1174]=12'b110001001010;
mem[1175]=12'b010011100110;
mem[1176]=12'b011110000011;
mem[1177]=12'b011100000100;
mem[1178]=12'b100101101110;
mem[1179]=12'b011111101000;
mem[1180]=12'b011100110110;
mem[1181]=12'b100001011011;
mem[1182]=12'b010110110011;
mem[1183]=12'b100001011001;
mem[1184]=12'b100000110010;
mem[1185]=12'b011111011111;
mem[1186]=12'b011101100011;
mem[1187]=12'b001010111101;
mem[1188]=12'b100000110101;
mem[1189]=12'b011111111111;
mem[1190]=12'b100011101110;
mem[1191]=12'b100010111001;
mem[1192]=12'b100110000011;
mem[1193]=12'b100011101100;
mem[1194]=12'b010101000100;
mem[1195]=12'b100011011111;
mem[1196]=12'b100011101011;
mem[1197]=12'b100100001000;
mem[1198]=12'b101100111100;
mem[1199]=12'b100001110110;
mem[1200]=12'b011001110101;
mem[1201]=12'b010110110001;
mem[1202]=12'b011101100110;
mem[1203]=12'b011000110001;
mem[1204]=12'b100010000011;
mem[1205]=12'b100010010100;
mem[1206]=12'b010100111001;
mem[1207]=12'b011110100011;
mem[1208]=12'b100010111011;
mem[1209]=12'b011110101011;
mem[1210]=12'b010110100101;
mem[1211]=12'b100010010000;
mem[1212]=12'b011000111000;
mem[1213]=12'b100001110000;
mem[1214]=12'b101011110101;
mem[1215]=12'b000100011111;
mem[1216]=12'b100000111110;
mem[1217]=12'b011111010101;
mem[1218]=12'b011000011111;
mem[1219]=12'b100010101100;
mem[1220]=12'b100000100000;
mem[1221]=12'b100000110100;
mem[1222]=12'b011011110010;
mem[1223]=12'b100010010011;
mem[1224]=12'b100001000011;
mem[1225]=12'b100111001000;
mem[1226]=12'b100000011110;
mem[1227]=12'b010001001101;
mem[1228]=12'b101011001000;
mem[1229]=12'b001110001010;
mem[1230]=12'b011101000010;
mem[1231]=12'b100001100101;
mem[1232]=12'b011001000011;
mem[1233]=12'b011111111100;
mem[1234]=12'b100000010011;
mem[1235]=12'b011110111111;
mem[1236]=12'b010000001010;
mem[1237]=12'b011111010110;
mem[1238]=12'b001110001101;
mem[1239]=12'b011111100100;
mem[1240]=12'b010111111100;
mem[1241]=12'b100101001111;
mem[1242]=12'b100001011010;
mem[1243]=12'b100001011110;
mem[1244]=12'b011110001110;
mem[1245]=12'b011011001001;
mem[1246]=12'b100011110110;
mem[1247]=12'b100111010001;
mem[1248]=12'b011100111001;
mem[1249]=12'b100001111000;
mem[1250]=12'b100001100110;
mem[1251]=12'b011010000001;
mem[1252]=12'b011111111111;
mem[1253]=12'b100101001101;
mem[1254]=12'b100011101010;
mem[1255]=12'b010100100011;
mem[1256]=12'b011101000101;
mem[1257]=12'b100000111110;
mem[1258]=12'b010111111011;
mem[1259]=12'b100110000000;
mem[1260]=12'b011010100001;
mem[1261]=12'b100011010010;
mem[1262]=12'b011101111101;
mem[1263]=12'b100001011101;
mem[1264]=12'b010111010000;
mem[1265]=12'b001110001001;
mem[1266]=12'b100100111110;
mem[1267]=12'b011000000010;
mem[1268]=12'b100011111000;
mem[1269]=12'b100011010100;
mem[1270]=12'b100101110000;
mem[1271]=12'b010100001100;
mem[1272]=12'b100101011011;
mem[1273]=12'b100011000110;
mem[1274]=12'b011000010001;
mem[1275]=12'b011101010010;
mem[1276]=12'b100100000001;
mem[1277]=12'b100010100000;
mem[1278]=12'b011110000110;
mem[1279]=12'b100001001110;
mem[1280]=12'b010110011000;
mem[1281]=12'b101001000000;
mem[1282]=12'b100001101111;
mem[1283]=12'b110101110111;
mem[1284]=12'b011011100111;
mem[1285]=12'b100010011100;
mem[1286]=12'b011110010100;
mem[1287]=12'b010101000000;
mem[1288]=12'b100001000110;
mem[1289]=12'b101010110011;
mem[1290]=12'b011110001001;
mem[1291]=12'b011001111110;
mem[1292]=12'b101010110011;
mem[1293]=12'b100010001101;
mem[1294]=12'b001010011110;
mem[1295]=12'b100100000011;
mem[1296]=12'b011110000101;
mem[1297]=12'b011101000010;
mem[1298]=12'b011100001111;
mem[1299]=12'b100010010010;
mem[1300]=12'b010111111011;
mem[1301]=12'b100001001101;
mem[1302]=12'b100011010000;
mem[1303]=12'b100001010000;
mem[1304]=12'b011101001000;
mem[1305]=12'b100011001011;
mem[1306]=12'b100011000100;
mem[1307]=12'b100001001001;
mem[1308]=12'b100100111100;
mem[1309]=12'b100010111100;
mem[1310]=12'b100001111000;
mem[1311]=12'b100111001011;
mem[1312]=12'b100001001100;
mem[1313]=12'b100011101011;
mem[1314]=12'b100000010000;
mem[1315]=12'b010000001010;
mem[1316]=12'b100010101101;
mem[1317]=12'b100001010111;
mem[1318]=12'b011011000111;
mem[1319]=12'b101010011001;
mem[1320]=12'b011001110110;
mem[1321]=12'b011110101100;
mem[1322]=12'b100010011000;
mem[1323]=12'b100100110111;
mem[1324]=12'b010110110000;
mem[1325]=12'b011110010010;
mem[1326]=12'b101101010000;
mem[1327]=12'b010001110011;
mem[1328]=12'b100000011001;
mem[1329]=12'b011111100101;
mem[1330]=12'b010101110011;
mem[1331]=12'b101010000110;
mem[1332]=12'b100000001101;
mem[1333]=12'b011110000011;
mem[1334]=12'b100001001101;
mem[1335]=12'b011111100111;
mem[1336]=12'b011101001011;
mem[1337]=12'b010110010011;
mem[1338]=12'b100000001101;
mem[1339]=12'b011111011101;
mem[1340]=12'b100100011000;
mem[1341]=12'b100010001000;
mem[1342]=12'b011011101011;
mem[1343]=12'b100001010010;
mem[1344]=12'b011111110110;
mem[1345]=12'b101010101010;
mem[1346]=12'b011011001001;
mem[1347]=12'b100011100110;
mem[1348]=12'b011110100011;
mem[1349]=12'b010100010010;
mem[1350]=12'b101101001011;
mem[1351]=12'b100010000111;
mem[1352]=12'b101011100011;
mem[1353]=12'b100110001011;
mem[1354]=12'b010110010010;
mem[1355]=12'b100100011100;
mem[1356]=12'b100010110001;
mem[1357]=12'b100011000110;
mem[1358]=12'b100010101110;
mem[1359]=12'b100010101111;
mem[1360]=12'b100010100011;
mem[1361]=12'b100010110100;
mem[1362]=12'b100010100111;
mem[1363]=12'b011100101010;
mem[1364]=12'b100100111100;
mem[1365]=12'b100100011000;
mem[1366]=12'b100001010100;
mem[1367]=12'b100110010001;
mem[1368]=12'b010010110101;
mem[1369]=12'b100010011010;
mem[1370]=12'b100001011100;
mem[1371]=12'b011111010011;
mem[1372]=12'b100100011101;
mem[1373]=12'b100001011100;
mem[1374]=12'b011101110001;
mem[1375]=12'b010101000010;
mem[1376]=12'b100000001110;
mem[1377]=12'b011111010010;
mem[1378]=12'b011000111011;
mem[1379]=12'b011011111110;
mem[1380]=12'b100000101000;
mem[1381]=12'b100001100100;
mem[1382]=12'b011001000010;
mem[1383]=12'b011001001110;
mem[1384]=12'b100000010011;
mem[1385]=12'b011111001011;
mem[1386]=12'b100111111111;
mem[1387]=12'b001100110011;
mem[1388]=12'b100001111011;
mem[1389]=12'b100100001011;
mem[1390]=12'b100000000010;
mem[1391]=12'b100000010010;
mem[1392]=12'b011110011011;
mem[1393]=12'b011001101000;
mem[1394]=12'b011111110001;
mem[1395]=12'b100001011001;
mem[1396]=12'b100010011011;
mem[1397]=12'b011111001101;
mem[1398]=12'b010111011111;
mem[1399]=12'b011101010011;
mem[1400]=12'b100000111001;
mem[1401]=12'b011101110110;
mem[1402]=12'b100000111011;
mem[1403]=12'b011100001111;
mem[1404]=12'b100111011110;
mem[1405]=12'b011111110101;
mem[1406]=12'b011000111110;
mem[1407]=12'b100101000011;
mem[1408]=12'b100000010101;
mem[1409]=12'b011011101101;
mem[1410]=12'b101010110100;
mem[1411]=12'b010101100111;
mem[1412]=12'b100010001111;
mem[1413]=12'b100001011101;
mem[1414]=12'b011011001110;
mem[1415]=12'b100010011011;
mem[1416]=12'b011110001110;
mem[1417]=12'b100011100000;
mem[1418]=12'b011011000111;
mem[1419]=12'b011111110011;
mem[1420]=12'b001010010101;
mem[1421]=12'b011011000001;
mem[1422]=12'b100110100100;
mem[1423]=12'b011100010011;
mem[1424]=12'b101010101001;
mem[1425]=12'b100011010111;
mem[1426]=12'b010101001000;
mem[1427]=12'b100001000111;
mem[1428]=12'b100001111101;
mem[1429]=12'b011110111101;
mem[1430]=12'b100001000101;
mem[1431]=12'b100001000011;
mem[1432]=12'b010111101111;
mem[1433]=12'b110011100010;
mem[1434]=12'b011101110011;
mem[1435]=12'b100001101001;
mem[1436]=12'b011000100100;
mem[1437]=12'b100111100110;
mem[1438]=12'b011111111011;
mem[1439]=12'b010111001111;
mem[1440]=12'b100100111101;
mem[1441]=12'b100101011111;
mem[1442]=12'b100000001001;
mem[1443]=12'b011111000100;
mem[1444]=12'b010111011111;
mem[1445]=12'b011111111101;
mem[1446]=12'b101000000010;
mem[1447]=12'b100001110011;
mem[1448]=12'b100011100001;
mem[1449]=12'b010000101110;
mem[1450]=12'b100000000111;
mem[1451]=12'b100100001111;
mem[1452]=12'b100011100010;
mem[1453]=12'b100000111101;
mem[1454]=12'b011100011101;
mem[1455]=12'b100011000111;
mem[1456]=12'b100000110100;
mem[1457]=12'b100111000011;
mem[1458]=12'b011010010110;
mem[1459]=12'b101000000000;
mem[1460]=12'b010111001110;
mem[1461]=12'b101011000111;
mem[1462]=12'b100001110100;
mem[1463]=12'b100101110000;
mem[1464]=12'b100110111011;
mem[1465]=12'b100001001010;
mem[1466]=12'b011010001010;
mem[1467]=12'b011101000010;
mem[1468]=12'b011010110101;
mem[1469]=12'b100100100001;
mem[1470]=12'b100101101111;
mem[1471]=12'b010101011111;
mem[1472]=12'b001000100111;
mem[1473]=12'b000000000011;
mem[1474]=12'b101100110111;
mem[1475]=12'b010101000000;
mem[1476]=12'b011101001101;
mem[1477]=12'b011010010000;
mem[1478]=12'b100010101000;
mem[1479]=12'b010110000000;
mem[1480]=12'b011100100001;
mem[1481]=12'b011011111010;
mem[1482]=12'b101010000101;
mem[1483]=12'b100000111000;
mem[1484]=12'b011111101000;
mem[1485]=12'b100000110000;
mem[1486]=12'b010000001000;
mem[1487]=12'b011111100010;
mem[1488]=12'b010111100011;
mem[1489]=12'b011011111011;
mem[1490]=12'b011101010110;
mem[1491]=12'b011111011111;
mem[1492]=12'b011111111001;
mem[1493]=12'b100011001000;
mem[1494]=12'b100000000001;
mem[1495]=12'b011110001101;
mem[1496]=12'b011111110000;
mem[1497]=12'b001011001001;
mem[1498]=12'b011110100010;
mem[1499]=12'b100001110111;
mem[1500]=12'b011001100111;
mem[1501]=12'b101110001010;
mem[1502]=12'b100011011100;
mem[1503]=12'b011010101001;
mem[1504]=12'b011101001100;
mem[1505]=12'b100001110010;
mem[1506]=12'b100001101000;
mem[1507]=12'b011111101100;
mem[1508]=12'b100011110001;
mem[1509]=12'b011100010100;
mem[1510]=12'b100001101011;
mem[1511]=12'b011111111111;
mem[1512]=12'b011110110010;
mem[1513]=12'b100001001000;
mem[1514]=12'b100010101010;
mem[1515]=12'b011111010100;
mem[1516]=12'b011101010011;
mem[1517]=12'b010101110000;
mem[1518]=12'b100000000000;
mem[1519]=12'b101010001110;
mem[1520]=12'b011111111110;
mem[1521]=12'b100011001110;
mem[1522]=12'b100001100010;
mem[1523]=12'b011111110101;
mem[1524]=12'b100101101000;
mem[1525]=12'b011110000111;
mem[1526]=12'b011000000010;
mem[1527]=12'b100101000011;
mem[1528]=12'b011001010111;
mem[1529]=12'b100110001010;
mem[1530]=12'b011100101010;
mem[1531]=12'b010110111001;
mem[1532]=12'b010011100001;
mem[1533]=12'b100010001101;
mem[1534]=12'b100011001110;
mem[1535]=12'b010110001111;
mem[1536]=12'b100111110011;
mem[1537]=12'b100001110001;
mem[1538]=12'b010111101011;
mem[1539]=12'b100000100101;
mem[1540]=12'b100010110000;
mem[1541]=12'b100001011010;
mem[1542]=12'b011110000101;
mem[1543]=12'b100000111001;
mem[1544]=12'b011110110100;
mem[1545]=12'b100000001010;
mem[1546]=12'b101011111100;
mem[1547]=12'b010101011100;
mem[1548]=12'b100001100000;
mem[1549]=12'b101011000001;
mem[1550]=12'b010001011011;
mem[1551]=12'b010010100110;
mem[1552]=12'b101000111011;
mem[1553]=12'b010111011001;
mem[1554]=12'b011110011111;
mem[1555]=12'b100000001100;
mem[1556]=12'b100001001010;
mem[1557]=12'b011110000011;
mem[1558]=12'b011011010100;
mem[1559]=12'b011101010000;
mem[1560]=12'b010101000001;
mem[1561]=12'b011010101111;
mem[1562]=12'b100001111011;
mem[1563]=12'b100001011010;
mem[1564]=12'b011010011010;
mem[1565]=12'b011111111101;
mem[1566]=12'b011111100010;
mem[1567]=12'b001101000011;
mem[1568]=12'b100100100111;
mem[1569]=12'b001011100010;
mem[1570]=12'b011111010110;
mem[1571]=12'b100010011101;
mem[1572]=12'b100100110111;
mem[1573]=12'b011010001110;
mem[1574]=12'b100000010101;
mem[1575]=12'b100110100110;
mem[1576]=12'b100010101010;
mem[1577]=12'b010111101100;
mem[1578]=12'b011111000111;
mem[1579]=12'b100000100100;
mem[1580]=12'b100111001011;
mem[1581]=12'b101001111101;
mem[1582]=12'b001010110100;
mem[1583]=12'b010111110101;
mem[1584]=12'b011111111010;
mem[1585]=12'b011100100100;
mem[1586]=12'b010110001110;
mem[1587]=12'b100000000001;
mem[1588]=12'b011101011000;
mem[1589]=12'b011100110010;
mem[1590]=12'b011011001000;
mem[1591]=12'b100001101001;
mem[1592]=12'b100011000100;
mem[1593]=12'b011101111010;
mem[1594]=12'b100011101010;
mem[1595]=12'b011010000100;
mem[1596]=12'b100101101011;
mem[1597]=12'b011100101101;
mem[1598]=12'b010010100011;
mem[1599]=12'b100001010001;
mem[1600]=12'b011111100010;
mem[1601]=12'b100000000101;
mem[1602]=12'b100011111100;
mem[1603]=12'b011000000110;
mem[1604]=12'b011111001100;
mem[1605]=12'b101010110100;
mem[1606]=12'b010001011111;
mem[1607]=12'b001011011001;
mem[1608]=12'b010100100010;
mem[1609]=12'b100001111101;
mem[1610]=12'b100001000000;
mem[1611]=12'b100110111000;
mem[1612]=12'b100001011101;
mem[1613]=12'b100001011000;
mem[1614]=12'b011011111011;
mem[1615]=12'b011110101001;
mem[1616]=12'b100010011001;
mem[1617]=12'b011011111100;
mem[1618]=12'b100101011000;
mem[1619]=12'b011110001101;
mem[1620]=12'b011011111000;
mem[1621]=12'b011111111100;
mem[1622]=12'b011111100010;
mem[1623]=12'b100001100100;
mem[1624]=12'b100101000101;
mem[1625]=12'b011101000101;
mem[1626]=12'b100011011111;
mem[1627]=12'b011000001100;
mem[1628]=12'b011110111101;
mem[1629]=12'b011010101001;
mem[1630]=12'b100001111111;
mem[1631]=12'b101001011000;
mem[1632]=12'b001110000000;
mem[1633]=12'b011111101111;
mem[1634]=12'b011110000011;
mem[1635]=12'b100001011000;
mem[1636]=12'b011110110001;
mem[1637]=12'b100001011101;
mem[1638]=12'b100100111001;
mem[1639]=12'b100001100111;
mem[1640]=12'b001011010000;
mem[1641]=12'b011110000011;
mem[1642]=12'b010101100100;
mem[1643]=12'b011110000010;
mem[1644]=12'b010001110000;
mem[1645]=12'b100001001110;
mem[1646]=12'b100111100010;
mem[1647]=12'b010111100101;
mem[1648]=12'b011110111100;
mem[1649]=12'b100100101000;
mem[1650]=12'b100001100011;
mem[1651]=12'b011111110011;
mem[1652]=12'b011100001000;
mem[1653]=12'b100001101110;
mem[1654]=12'b100000000111;
mem[1655]=12'b101010110111;
mem[1656]=12'b100010000100;
mem[1657]=12'b100010110100;
mem[1658]=12'b100011011110;
mem[1659]=12'b100010101110;
mem[1660]=12'b010110101110;
mem[1661]=12'b011101101000;
mem[1662]=12'b100011011010;
mem[1663]=12'b100010000100;
mem[1664]=12'b100010100111;
mem[1665]=12'b100100000001;
mem[1666]=12'b010001010011;
mem[1667]=12'b011111111000;
mem[1668]=12'b100000000111;
mem[1669]=12'b100001001011;
mem[1670]=12'b100100001110;
mem[1671]=12'b011001010100;
mem[1672]=12'b100000000010;
mem[1673]=12'b100001011101;
mem[1674]=12'b100110000000;
mem[1675]=12'b001010011101;
mem[1676]=12'b011111101000;
mem[1677]=12'b100010000110;
mem[1678]=12'b011111011001;
mem[1679]=12'b100000111000;
mem[1680]=12'b100000010100;
mem[1681]=12'b101000110100;
mem[1682]=12'b011010100100;
mem[1683]=12'b100000111101;
mem[1684]=12'b011110110010;
mem[1685]=12'b011111111100;
mem[1686]=12'b011111010110;
mem[1687]=12'b100010100000;
mem[1688]=12'b011000000111;
mem[1689]=12'b011110011000;
mem[1690]=12'b100010101111;
mem[1691]=12'b011101100011;
mem[1692]=12'b011111010000;
mem[1693]=12'b011001101101;
mem[1694]=12'b010001001100;
mem[1695]=12'b011111110111;
mem[1696]=12'b100011011110;
mem[1697]=12'b011110001001;
mem[1698]=12'b100001111101;
mem[1699]=12'b011001111011;
mem[1700]=12'b011110101001;
mem[1701]=12'b011001101011;
mem[1702]=12'b100000000100;
mem[1703]=12'b011110100011;
mem[1704]=12'b100001001010;
mem[1705]=12'b011010001110;
mem[1706]=12'b100010111111;
mem[1707]=12'b011110100111;
mem[1708]=12'b100001100010;
mem[1709]=12'b100000101110;
mem[1710]=12'b100010110001;
mem[1711]=12'b101001000110;
mem[1712]=12'b101011001110;
mem[1713]=12'b010101111010;
mem[1714]=12'b100010100011;
mem[1715]=12'b010010110010;
mem[1716]=12'b100010001100;
mem[1717]=12'b100000110110;
mem[1718]=12'b100011100101;
mem[1719]=12'b100010100101;
mem[1720]=12'b100011001110;
mem[1721]=12'b100010010111;
mem[1722]=12'b100001100001;
mem[1723]=12'b011011000001;
mem[1724]=12'b011110010010;
mem[1725]=12'b100010110001;
mem[1726]=12'b100110100100;
mem[1727]=12'b100001010111;
mem[1728]=12'b011110011001;
mem[1729]=12'b011000100110;
mem[1730]=12'b010110000100;
mem[1731]=12'b100111101001;
mem[1732]=12'b100010000110;
mem[1733]=12'b100001110000;
mem[1734]=12'b011111111101;
mem[1735]=12'b010001101101;
mem[1736]=12'b100001110000;
mem[1737]=12'b100110011010;
mem[1738]=12'b100001100000;
mem[1739]=12'b011001110100;
mem[1740]=12'b011101010000;
mem[1741]=12'b100110100111;
mem[1742]=12'b100010011000;
mem[1743]=12'b101001001100;
mem[1744]=12'b100010000000;
mem[1745]=12'b101101101000;
mem[1746]=12'b100010010111;
mem[1747]=12'b100011010010;
mem[1748]=12'b100110001100;
mem[1749]=12'b010011010100;
mem[1750]=12'b011100100111;
mem[1751]=12'b011111111011;
mem[1752]=12'b100000000111;
mem[1753]=12'b001001011111;
mem[1754]=12'b100110000110;
mem[1755]=12'b100001010000;
mem[1756]=12'b011111010000;
mem[1757]=12'b100011101101;
mem[1758]=12'b100010100010;
mem[1759]=12'b011101000000;
mem[1760]=12'b011011000110;
mem[1761]=12'b011111101110;
mem[1762]=12'b101101110010;
mem[1763]=12'b100001001111;
mem[1764]=12'b100110110100;
mem[1765]=12'b100000011000;
mem[1766]=12'b100001010011;
mem[1767]=12'b101010011010;
mem[1768]=12'b010110011110;
mem[1769]=12'b011100111111;
mem[1770]=12'b100010000000;
mem[1771]=12'b011011101110;
mem[1772]=12'b011010000110;
mem[1773]=12'b100100000111;
mem[1774]=12'b100001110010;
mem[1775]=12'b011100001101;
mem[1776]=12'b001111110001;
mem[1777]=12'b100000111001;
mem[1778]=12'b100110001111;
mem[1779]=12'b011110100001;
mem[1780]=12'b100001100111;
mem[1781]=12'b010111001110;
mem[1782]=12'b011011101111;
mem[1783]=12'b101000100001;
mem[1784]=12'b011100111111;
mem[1785]=12'b100001101001;
mem[1786]=12'b011101001100;
mem[1787]=12'b100100101101;
mem[1788]=12'b011101010000;
mem[1789]=12'b100001011010;
mem[1790]=12'b100001100011;
mem[1791]=12'b100101110000;
mem[1792]=12'b010010010001;
mem[1793]=12'b100011001111;
mem[1794]=12'b100001001101;
mem[1795]=12'b100000010000;
mem[1796]=12'b011111000010;
mem[1797]=12'b100000001101;
mem[1798]=12'b100101010101;
mem[1799]=12'b011000111011;
mem[1800]=12'b100001010101;
mem[1801]=12'b011101101101;
mem[1802]=12'b011100001000;
mem[1803]=12'b011101111101;
mem[1804]=12'b011001101100;
mem[1805]=12'b100010111001;
mem[1806]=12'b011111001000;
mem[1807]=12'b100001100101;
mem[1808]=12'b010111100100;
mem[1809]=12'b011111110000;
mem[1810]=12'b011111001011;
mem[1811]=12'b011111101011;
mem[1812]=12'b100010010001;
mem[1813]=12'b011101101100;
mem[1814]=12'b011101101111;
mem[1815]=12'b100000110101;
mem[1816]=12'b100100010000;
mem[1817]=12'b011110001011;
mem[1818]=12'b010011011011;
mem[1819]=12'b011010010010;
mem[1820]=12'b011111101111;
mem[1821]=12'b100000111001;
mem[1822]=12'b100111110100;
mem[1823]=12'b001000011101;
mem[1824]=12'b100000000011;
mem[1825]=12'b100000110101;
mem[1826]=12'b011111011111;
mem[1827]=12'b001011111001;
mem[1828]=12'b100011010101;
mem[1829]=12'b011000101011;
mem[1830]=12'b100010110001;
mem[1831]=12'b101011110001;
mem[1832]=12'b100001111101;
mem[1833]=12'b011100000001;
mem[1834]=12'b000100010011;
mem[1835]=12'b100001101000;
mem[1836]=12'b011100011010;
mem[1837]=12'b100010100011;
mem[1838]=12'b100000001100;
mem[1839]=12'b001000111100;
mem[1840]=12'b011111110001;
mem[1841]=12'b011111101010;
mem[1842]=12'b100001010101;
mem[1843]=12'b100010101110;
mem[1844]=12'b100001001101;
mem[1845]=12'b011110011010;
mem[1846]=12'b101000010111;
mem[1847]=12'b100000001011;
mem[1848]=12'b011000100001;
mem[1849]=12'b011111110011;
mem[1850]=12'b101100010101;
mem[1851]=12'b001001011100;
mem[1852]=12'b011110111000;
mem[1853]=12'b011010011011;
mem[1854]=12'b011000000111;
mem[1855]=12'b011101101011;
mem[1856]=12'b100010001010;
mem[1857]=12'b100101110000;
mem[1858]=12'b011011110011;
mem[1859]=12'b011001111011;
mem[1860]=12'b100011100000;
mem[1861]=12'b011101111001;
mem[1862]=12'b100000000111;
mem[1863]=12'b100010010100;
mem[1864]=12'b100100101011;
mem[1865]=12'b010111010000;
mem[1866]=12'b011101011001;
mem[1867]=12'b011011110001;
mem[1868]=12'b100010110010;
mem[1869]=12'b100001001000;
mem[1870]=12'b100100000011;
mem[1871]=12'b011110101110;
mem[1872]=12'b100001001010;
mem[1873]=12'b011111100101;
mem[1874]=12'b100010000000;
mem[1875]=12'b100101101111;
mem[1876]=12'b100000000110;
mem[1877]=12'b011010011010;
mem[1878]=12'b100101101101;
mem[1879]=12'b100001001101;
mem[1880]=12'b011111111010;
mem[1881]=12'b011111101101;
mem[1882]=12'b100000000100;
mem[1883]=12'b011011000011;
mem[1884]=12'b100101001111;
mem[1885]=12'b011100110111;
mem[1886]=12'b100001000001;
mem[1887]=12'b011110010011;
mem[1888]=12'b010101011110;
mem[1889]=12'b011011010010;
mem[1890]=12'b100101000010;
mem[1891]=12'b101010101111;
mem[1892]=12'b011011100110;
mem[1893]=12'b001100000101;
mem[1894]=12'b100101001101;
mem[1895]=12'b011010011100;
mem[1896]=12'b011110101110;
mem[1897]=12'b100110101010;
mem[1898]=12'b010011100010;
mem[1899]=12'b011010101111;
mem[1900]=12'b011110110011;
mem[1901]=12'b011111110100;
mem[1902]=12'b100001010111;
mem[1903]=12'b101100000110;
mem[1904]=12'b011011110000;
mem[1905]=12'b110010001100;
mem[1906]=12'b100010010000;
mem[1907]=12'b101001001000;
mem[1908]=12'b100001000111;
mem[1909]=12'b011101101000;
mem[1910]=12'b010100100100;
mem[1911]=12'b100000111010;
mem[1912]=12'b101000011000;
mem[1913]=12'b010111110101;
mem[1914]=12'b011111010001;
mem[1915]=12'b100000000001;
mem[1916]=12'b100100010100;
mem[1917]=12'b001011010111;
mem[1918]=12'b100011001001;
mem[1919]=12'b010001110111;
mem[1920]=12'b011111110100;
mem[1921]=12'b011000001010;
mem[1922]=12'b011001101101;
mem[1923]=12'b100100110001;
mem[1924]=12'b100011011100;
mem[1925]=12'b100010011100;
mem[1926]=12'b100011110001;
mem[1927]=12'b011001101110;
mem[1928]=12'b010101001110;
mem[1929]=12'b100001111110;
mem[1930]=12'b101001010011;
mem[1931]=12'b100010010111;
mem[1932]=12'b011000011011;
mem[1933]=12'b100010011100;
mem[1934]=12'b100011011111;
mem[1935]=12'b010001001001;
mem[1936]=12'b100001010100;
mem[1937]=12'b010010010100;
mem[1938]=12'b100001010010;
mem[1939]=12'b011001010101;
mem[1940]=12'b100001011000;
mem[1941]=12'b011101010101;
mem[1942]=12'b100010011101;
mem[1943]=12'b100001111000;
mem[1944]=12'b100000011100;
mem[1945]=12'b101011000011;
mem[1946]=12'b100011100101;
mem[1947]=12'b100001111110;
mem[1948]=12'b011101101100;
mem[1949]=12'b010100000110;
mem[1950]=12'b100010001001;
mem[1951]=12'b101010010000;
mem[1952]=12'b011100110011;
mem[1953]=12'b010111000010;
mem[1954]=12'b011111111110;
mem[1955]=12'b011101111110;
mem[1956]=12'b001100000011;
mem[1957]=12'b011110101101;
mem[1958]=12'b010110011010;
mem[1959]=12'b011010010110;
mem[1960]=12'b100010100011;
mem[1961]=12'b100001001001;
mem[1962]=12'b001110110101;
mem[1963]=12'b011101101110;
mem[1964]=12'b011100100110;
mem[1965]=12'b011111100001;
mem[1966]=12'b011001000010;
mem[1967]=12'b100011001101;
mem[1968]=12'b011110000100;
mem[1969]=12'b100011000100;
mem[1970]=12'b100000010111;
mem[1971]=12'b101000111100;
mem[1972]=12'b100111110100;
mem[1973]=12'b100001011010;
mem[1974]=12'b011111100110;
mem[1975]=12'b011010010110;
mem[1976]=12'b011101110110;
mem[1977]=12'b100001100110;
mem[1978]=12'b100000100011;
mem[1979]=12'b100111101100;
mem[1980]=12'b100000000100;
mem[1981]=12'b100100000001;
mem[1982]=12'b011110000011;
mem[1983]=12'b100001110101;
mem[1984]=12'b100000011110;
mem[1985]=12'b011100101110;
mem[1986]=12'b100001100100;
mem[1987]=12'b011111011001;
mem[1988]=12'b101001100101;
mem[1989]=12'b100001011101;
mem[1990]=12'b011000110100;
mem[1991]=12'b100000001001;
mem[1992]=12'b100011001010;
mem[1993]=12'b011111000110;
mem[1994]=12'b011100001001;
mem[1995]=12'b011101011110;
mem[1996]=12'b010010110100;
mem[1997]=12'b100001011001;
mem[1998]=12'b100011001001;
mem[1999]=12'b011010000111;
mem[2000]=12'b100001100001;
mem[2001]=12'b011111011010;
mem[2002]=12'b100001101000;
mem[2003]=12'b101110110011;
mem[2004]=12'b011101011010;
mem[2005]=12'b100001111110;
mem[2006]=12'b011100111011;
mem[2007]=12'b100010010011;
mem[2008]=12'b100010110000;
mem[2009]=12'b100000111011;
mem[2010]=12'b001100000011;
mem[2011]=12'b100111000000;
mem[2012]=12'b011110000001;
mem[2013]=12'b011001111001;
mem[2014]=12'b100001100111;
mem[2015]=12'b100100011010;
mem[2016]=12'b001011001000;
mem[2017]=12'b011011110111;
mem[2018]=12'b011011110100;
mem[2019]=12'b100001000001;
mem[2020]=12'b101110101011;
mem[2021]=12'b100100000011;
mem[2022]=12'b100001001110;
mem[2023]=12'b100010101011;
mem[2024]=12'b100001100011;
mem[2025]=12'b101000111000;
mem[2026]=12'b010010110111;
mem[2027]=12'b101000011000;
mem[2028]=12'b011011011011;
mem[2029]=12'b100110000001;
mem[2030]=12'b100101011101;
mem[2031]=12'b100101011011;
mem[2032]=12'b100001011101;
mem[2033]=12'b011111010110;
mem[2034]=12'b100011000000;
mem[2035]=12'b011000100110;
mem[2036]=12'b010010000110;
mem[2037]=12'b100000111100;
mem[2038]=12'b101100111101;
mem[2039]=12'b011101110011;
mem[2040]=12'b100001001101;
mem[2041]=12'b100001000010;
mem[2042]=12'b011110000011;
mem[2043]=12'b011100010100;
mem[2044]=12'b011011000001;
mem[2045]=12'b100001001001;
mem[2046]=12'b110000101100;
mem[2047]=12'b011101111001;
mem[2048]=12'b001001011011;
mem[2049]=12'b100000000110;
mem[2050]=12'b100100011000;
mem[2051]=12'b100000111000;
mem[2052]=12'b011000010010;
mem[2053]=12'b101010000111;
mem[2054]=12'b011001101110;
mem[2055]=12'b100110000110;
mem[2056]=12'b100001000111;
mem[2057]=12'b100000010111;
mem[2058]=12'b110011100000;
mem[2059]=12'b100100100110;
mem[2060]=12'b011111101001;
mem[2061]=12'b000111010100;
mem[2062]=12'b100100011110;
mem[2063]=12'b011010111111;
mem[2064]=12'b011101101011;
mem[2065]=12'b011100000010;
mem[2066]=12'b100001001010;
mem[2067]=12'b100000100100;
mem[2068]=12'b100000011000;
mem[2069]=12'b100101000100;
mem[2070]=12'b100010011011;
mem[2071]=12'b001010110010;
mem[2072]=12'b101011000110;
mem[2073]=12'b011110100100;
mem[2074]=12'b001110110110;
mem[2075]=12'b100001101011;
mem[2076]=12'b010110110010;
mem[2077]=12'b100011111101;
mem[2078]=12'b101011011010;
mem[2079]=12'b011011011101;
mem[2080]=12'b100011011100;
mem[2081]=12'b100010110001;
mem[2082]=12'b101001101001;
mem[2083]=12'b100001000010;
mem[2084]=12'b011011100000;
mem[2085]=12'b100011101110;
mem[2086]=12'b000100101110;
mem[2087]=12'b011111110110;
mem[2088]=12'b100011000011;
mem[2089]=12'b100010000000;
mem[2090]=12'b100010001100;
mem[2091]=12'b100001010011;
mem[2092]=12'b011010100100;
mem[2093]=12'b100000000111;
mem[2094]=12'b010110011001;
mem[2095]=12'b101100100110;
mem[2096]=12'b100000010100;
mem[2097]=12'b101110110110;
mem[2098]=12'b100001000001;
mem[2099]=12'b011111101011;
mem[2100]=12'b011101000111;
mem[2101]=12'b100010110101;
mem[2102]=12'b011000111000;
mem[2103]=12'b011111110100;
mem[2104]=12'b100000000000;
mem[2105]=12'b100011100101;
mem[2106]=12'b011101101110;
mem[2107]=12'b100001001111;
mem[2108]=12'b010110001000;
mem[2109]=12'b100101100100;
mem[2110]=12'b100010011001;
mem[2111]=12'b011101101100;
mem[2112]=12'b101011010101;
mem[2113]=12'b100010101111;
mem[2114]=12'b011101111110;
mem[2115]=12'b011100010100;
mem[2116]=12'b100001001100;
mem[2117]=12'b100100111011;
mem[2118]=12'b100011110110;
mem[2119]=12'b011001000011;
mem[2120]=12'b100100001000;
mem[2121]=12'b011110000010;
mem[2122]=12'b011000000101;
mem[2123]=12'b100111010111;
mem[2124]=12'b011100000110;
mem[2125]=12'b001101001101;
mem[2126]=12'b100000111000;
mem[2127]=12'b100010101111;
mem[2128]=12'b011110100011;
mem[2129]=12'b010011011011;
mem[2130]=12'b011100100010;
mem[2131]=12'b100110100100;
mem[2132]=12'b100001001011;
mem[2133]=12'b011010110011;
mem[2134]=12'b101001101111;
end

always@(posedge clk)
begin
  if (we) begin
    mem[addr] <= din;
  end
end

always @(posedge clk) dout <= mem[addr];

endmodule
