`timescale 1ns/1ps
module STAGE_THRESHOLD_ROM(
  addr,
  clk,
  din,
  dout,
  we);

input [4 : 0] addr;
input clk;
input [18 : 0] din;
output reg [18 : 0] dout;
input we;

reg [18:0] mem [0:31];

initial begin
mem[0]=19'b0000000110100101001;
mem[1]=19'b0000110111101001110;
mem[2]=19'b0001001011111111010;
mem[3]=19'b0010010011010011011;
mem[4]=19'b0001111010100110000;
mem[5]=19'b0010101000000101011;
mem[6]=19'b0010111111010110011;
mem[7]=19'b0011000100001110010;
mem[8]=19'b0011011001001110100;
mem[9]=19'b0100010100011011101;
mem[10]=19'b0100111000110110111;
mem[11]=19'b0110010100111000101;
mem[12]=19'b0110110100111101011;
mem[13]=19'b0110010001010110111;
mem[14]=19'b1000010101010110100;
mem[15]=19'b1000011101100101111;
mem[16]=19'b1000101001110101101;
mem[17]=19'b1001111001111111100;
mem[18]=19'b1010111101100100010;
mem[19]=19'b1011010010000001101;
mem[20]=19'b1101000101111111100;
mem[21]=19'b1101001110000101101;
end

always@(posedge clk)
begin
  if (we) begin
    mem[addr] <= din;
  end
end

always @(posedge clk) dout <= mem[addr];

endmodule