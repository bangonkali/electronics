`timescale 1ns/1ps
module FEAT_THRESHOLD_ROM(
  addr,
  clk,
  din,
  dout,
  we);

input [11 : 0] addr;
input clk;
input [16 : 0] din;
output reg [16 : 0] dout;
input we;

reg [16:0] mem [0:4095];

initial begin
mem[0]=17'b00000000110011011;
mem[1]=17'b00000011000001111;
mem[2]=17'b00000000110101111;
mem[3]=17'b00000000010100110;
mem[4]=17'b00000000011101010;
mem[5]=17'b00000001000000000;
mem[6]=17'b00000001100101111;
mem[7]=17'b11111111010011000;
mem[8]=17'b00000111010101010;
mem[9]=17'b00000001110111100;
mem[10]=17'b00000001101111010;
mem[11]=17'b00000000001110101;
mem[12]=17'b11111111100100100;
mem[13]=17'b00000000011011001;
mem[14]=17'b11101101001101100;
mem[15]=17'b00000000010001101;
mem[16]=17'b00001110100111001;
mem[17]=17'b00000000000100101;
mem[18]=17'b11111110110010101;
mem[19]=17'b11111100101100110;
mem[20]=17'b00000000100010101;
mem[21]=17'b00000000100011111;
mem[22]=17'b11111111101100011;
mem[23]=17'b11111111111000111;
mem[24]=17'b00000000011000101;
mem[25]=17'b11111110111111110;
mem[26]=17'b00000000100001101;
mem[27]=17'b11111111101100110;
mem[28]=17'b11111101111110000;
mem[29]=17'b11111101100111000;
mem[30]=17'b00000000111110100;
mem[31]=17'b11101111111110011;
mem[32]=17'b00000000001101100;
mem[33]=17'b11111111101110111;
mem[34]=17'b11110101000101001;
mem[35]=17'b00000000100101001;
mem[36]=17'b00000000001001100;
mem[37]=17'b00000000110111000;
mem[38]=17'b00000000111001100;
mem[39]=17'b00000100110100111;
mem[40]=17'b00000000011000100;
mem[41]=17'b11111111111110011;
mem[42]=17'b00000000000110100;
mem[43]=17'b00000000110101100;
mem[44]=17'b00000001000001010;
mem[45]=17'b11111111100100101;
mem[46]=17'b11111111011011000;
mem[47]=17'b11111011101011100;
mem[48]=17'b11111111000100110;
mem[49]=17'b00000000000111100;
mem[50]=17'b00001010110001101;
mem[51]=17'b00000000011000001;
mem[52]=17'b11111111100001110;
mem[53]=17'b00000100110011011;
mem[54]=17'b00000000000010101;
mem[55]=17'b00000000001010110;
mem[56]=17'b00000000010010000;
mem[57]=17'b00000000010010101;
mem[58]=17'b00000000010100111;
mem[59]=17'b00000000001010101;
mem[60]=17'b11111111100101001;
mem[61]=17'b11111111110110101;
mem[62]=17'b00000000101001110;
mem[63]=17'b00000000001011011;
mem[64]=17'b11111100111100011;
mem[65]=17'b00000000111101111;
mem[66]=17'b11111111110100011;
mem[67]=17'b11111110110001101;
mem[68]=17'b11111111111010011;
mem[69]=17'b00000100100001111;
mem[70]=17'b11111111101000000;
mem[71]=17'b00000001011010101;
mem[72]=17'b00000000010110001;
mem[73]=17'b11111110101000011;
mem[74]=17'b11111111111111111;
mem[75]=17'b00000101111001010;
mem[76]=17'b00000001101000001;
mem[77]=17'b00000100001100000;
mem[78]=17'b11111110000101101;
mem[79]=17'b11111111111100100;
mem[80]=17'b00000000010101011;
mem[81]=17'b00000000001000111;
mem[82]=17'b00000000001010000;
mem[83]=17'b11111111011011100;
mem[84]=17'b11111111001111010;
mem[85]=17'b00000000010100010;
mem[86]=17'b00000010000001000;
mem[87]=17'b11110011010010111;
mem[88]=17'b11111110001011100;
mem[89]=17'b11111111100001010;
mem[90]=17'b00000000010011011;
mem[91]=17'b00000011100110010;
mem[92]=17'b11111110101101100;
mem[93]=17'b11111101101000000;
mem[94]=17'b00000000010000010;
mem[95]=17'b00000000001110100;
mem[96]=17'b11111111001001100;
mem[97]=17'b11111111011010001;
mem[98]=17'b11111110001110111;
mem[99]=17'b11111110101011000;
mem[100]=17'b00000000110011001;
mem[101]=17'b11111111001011010;
mem[102]=17'b00000011000111111;
mem[103]=17'b11111101111011100;
mem[104]=17'b11111110001111100;
mem[105]=17'b00100000011101000;
mem[106]=17'b00000000111010010;
mem[107]=17'b11111111100100110;
mem[108]=17'b11111101010111000;
mem[109]=17'b11110010110011010;
mem[110]=17'b00000001100101010;
mem[111]=17'b00000100001011011;
mem[112]=17'b00000000001111010;
mem[113]=17'b11111111101000001;
mem[114]=17'b11111111111101100;
mem[115]=17'b11111111110101110;
mem[116]=17'b11111111100000110;
mem[117]=17'b00000000000110011;
mem[118]=17'b00000000110011100;
mem[119]=17'b11111101000111001;
mem[120]=17'b00000000011010000;
mem[121]=17'b11111111101011011;
mem[122]=17'b00000000101010110;
mem[123]=17'b00000000010100111;
mem[124]=17'b00000110000011001;
mem[125]=17'b00000111011100110;
mem[126]=17'b11111010111110101;
mem[127]=17'b11111110111100001;
mem[128]=17'b00000000001111011;
mem[129]=17'b11111011100111101;
mem[130]=17'b00000001000101010;
mem[131]=17'b00001101111111010;
mem[132]=17'b00000000000100011;
mem[133]=17'b00000000010000001;
mem[134]=17'b00000100100010110;
mem[135]=17'b11111111101000111;
mem[136]=17'b00000000101010110;
mem[137]=17'b00000000000101001;
mem[138]=17'b00000010100011000;
mem[139]=17'b11111110100010100;
mem[140]=17'b11110100100111001;
mem[141]=17'b11111110111111111;
mem[142]=17'b00000001001101001;
mem[143]=17'b00000000110010011;
mem[144]=17'b11111111010001010;
mem[145]=17'b11111111001110111;
mem[146]=17'b11111110100100000;
mem[147]=17'b11110101011100010;
mem[148]=17'b11111110011010010;
mem[149]=17'b11111111011101000;
mem[150]=17'b11111111101000011;
mem[151]=17'b00000011001011110;
mem[152]=17'b11111111101111111;
mem[153]=17'b00000001010000011;
mem[154]=17'b11111110110000011;
mem[155]=17'b11111101100100110;
mem[156]=17'b11111111001101111;
mem[157]=17'b00000000010100011;
mem[158]=17'b00000011100011100;
mem[159]=17'b00000000001000010;
mem[160]=17'b11111111111100011;
mem[161]=17'b00000000010100100;
mem[162]=17'b11101100011100111;
mem[163]=17'b00000000000111000;
mem[164]=17'b11111101011011100;
mem[165]=17'b00000000110101001;
mem[166]=17'b00000000010101111;
mem[167]=17'b00000001100000010;
mem[168]=17'b00000000011100110;
mem[169]=17'b00001010011001101;
mem[170]=17'b00000010011010101;
mem[171]=17'b00000000000000001;
mem[172]=17'b00000000000000000;
mem[173]=17'b11111111000101001;
mem[174]=17'b00000000011001101;
mem[175]=17'b00000000111001101;
mem[176]=17'b00000010010110010;
mem[177]=17'b11110100010101101;
mem[178]=17'b00000000000011000;
mem[179]=17'b11111110011100000;
mem[180]=17'b11111101110100111;
mem[181]=17'b11111111011100100;
mem[182]=17'b11111111110110000;
mem[183]=17'b00000010110001100;
mem[184]=17'b11111011010001000;
mem[185]=17'b11111111111111111;
mem[186]=17'b00000000101110010;
mem[187]=17'b11111100000010011;
mem[188]=17'b11111111001111010;
mem[189]=17'b11111111000000011;
mem[190]=17'b00000000011100101;
mem[191]=17'b00000010011101001;
mem[192]=17'b11111111011011100;
mem[193]=17'b11111111001111101;
mem[194]=17'b11111111110000100;
mem[195]=17'b00000010000010000;
mem[196]=17'b11111100110001000;
mem[197]=17'b00000011110110111;
mem[198]=17'b11111111010110100;
mem[199]=17'b11111110001000000;
mem[200]=17'b11111101011110110;
mem[201]=17'b11111010111000001;
mem[202]=17'b11111111111111001;
mem[203]=17'b11101110001010001;
mem[204]=17'b11111111011100101;
mem[205]=17'b00000000000011011;
mem[206]=17'b00000000010010111;
mem[207]=17'b11111111101000001;
mem[208]=17'b11111111101010001;
mem[209]=17'b11111111100111111;
mem[210]=17'b11111110111100010;
mem[211]=17'b11110110101010110;
mem[212]=17'b11111111110101111;
mem[213]=17'b00000010111110100;
mem[214]=17'b11111111110000101;
mem[215]=17'b00000001001101100;
mem[216]=17'b11111111011111110;
mem[217]=17'b11111110110100100;
mem[218]=17'b00000001001000100;
mem[219]=17'b11111111011001010;
mem[220]=17'b00000000100110001;
mem[221]=17'b11110000110101010;
mem[222]=17'b00000011110110100;
mem[223]=17'b00000000000010011;
mem[224]=17'b00000101110111111;
mem[225]=17'b00000000001101010;
mem[226]=17'b00000000100001011;
mem[227]=17'b00000000001100011;
mem[228]=17'b00000000000111100;
mem[229]=17'b11101011101100000;
mem[230]=17'b00000111001110110;
mem[231]=17'b00000000101100010;
mem[232]=17'b00000011111010010;
mem[233]=17'b11111111100010100;
mem[234]=17'b11111111101000010;
mem[235]=17'b11111111110100000;
mem[236]=17'b11111110111101000;
mem[237]=17'b00000000000001100;
mem[238]=17'b00000000001111001;
mem[239]=17'b11111101110100110;
mem[240]=17'b00000000010110001;
mem[241]=17'b11111110101100110;
mem[242]=17'b11111111110000100;
mem[243]=17'b11111101111011100;
mem[244]=17'b00000000000111001;
mem[245]=17'b00000011000011110;
mem[246]=17'b11111011101011110;
mem[247]=17'b11100110010101010;
mem[248]=17'b11111111100010110;
mem[249]=17'b00001111111110111;
mem[250]=17'b11110000000111010;
mem[251]=17'b11111110111100100;
mem[252]=17'b00000000001101011;
mem[253]=17'b00000000000011010;
mem[254]=17'b11111111010001110;
mem[255]=17'b00000010010010001;
mem[256]=17'b11111111100110100;
mem[257]=17'b11111110000000100;
mem[258]=17'b00000000001001010;
mem[259]=17'b00000000001000001;
mem[260]=17'b00000000111010001;
mem[261]=17'b00000000000001001;
mem[262]=17'b11111110010001010;
mem[263]=17'b00000001100111000;
mem[264]=17'b00000000000101100;
mem[265]=17'b11111111111110110;
mem[266]=17'b11111111110001101;
mem[267]=17'b00000001010010011;
mem[268]=17'b11110100101000101;
mem[269]=17'b00000000110100000;
mem[270]=17'b00000000000000100;
mem[271]=17'b00000001001111000;
mem[272]=17'b00000001010011001;
mem[273]=17'b11111111110011000;
mem[274]=17'b11111110111010101;
mem[275]=17'b11111111110010100;
mem[276]=17'b00000000001000100;
mem[277]=17'b11111111111100100;
mem[278]=17'b00000000110110001;
mem[279]=17'b11111111010110000;
mem[280]=17'b00000000000001111;
mem[281]=17'b00000000000000000;
mem[282]=17'b11111101000011000;
mem[283]=17'b00000100111001011;
mem[284]=17'b11111111111011010;
mem[285]=17'b00000000000000000;
mem[286]=17'b11111100111110110;
mem[287]=17'b11111111001111000;
mem[288]=17'b00000011011000101;
mem[289]=17'b11111111011001000;
mem[290]=17'b00000000101001001;
mem[291]=17'b11111111001100111;
mem[292]=17'b00000001011110111;
mem[293]=17'b11111110001110100;
mem[294]=17'b00000000100010111;
mem[295]=17'b11111111100000000;
mem[296]=17'b11111110011001000;
mem[297]=17'b11111111110011100;
mem[298]=17'b11111110110100111;
mem[299]=17'b11111111000110100;
mem[300]=17'b11111110111010100;
mem[301]=17'b11111111110110100;
mem[302]=17'b00000000000000001;
mem[303]=17'b00001000001001101;
mem[304]=17'b00000001010101001;
mem[305]=17'b00000000111010100;
mem[306]=17'b00000001010011100;
mem[307]=17'b11111101010001010;
mem[308]=17'b00000101011110001;
mem[309]=17'b00000000000111111;
mem[310]=17'b11111111010101110;
mem[311]=17'b11111101111000000;
mem[312]=17'b00000011111000110;
mem[313]=17'b11111110111001101;
mem[314]=17'b00000000011001000;
mem[315]=17'b11111110001110010;
mem[316]=17'b00010000101110100;
mem[317]=17'b00000000001111101;
mem[318]=17'b00000001001001110;
mem[319]=17'b11111111101011000;
mem[320]=17'b00000000101011101;
mem[321]=17'b11111101110010011;
mem[322]=17'b00000110111110010;
mem[323]=17'b00000000001000011;
mem[324]=17'b11111011001000100;
mem[325]=17'b00000000000111100;
mem[326]=17'b00000000011101011;
mem[327]=17'b11111111001111101;
mem[328]=17'b11100101001010010;
mem[329]=17'b00000000001001101;
mem[330]=17'b11110111111001001;
mem[331]=17'b00000000010000000;
mem[332]=17'b11111110100001000;
mem[333]=17'b00000000000110100;
mem[334]=17'b11111111101111101;
mem[335]=17'b11111111101000101;
mem[336]=17'b00000101011111110;
mem[337]=17'b00000000011100101;
mem[338]=17'b11111110001110101;
mem[339]=17'b00000000110101011;
mem[340]=17'b11111111101010001;
mem[341]=17'b00000001010011100;
mem[342]=17'b11111110000110000;
mem[343]=17'b00000101000011111;
mem[344]=17'b00000111010010101;
mem[345]=17'b00000100001010111;
mem[346]=17'b11111111110100111;
mem[347]=17'b11111111111111111;
mem[348]=17'b11111111110101010;
mem[349]=17'b00000000101110001;
mem[350]=17'b11111110101001000;
mem[351]=17'b11110110100110001;
mem[352]=17'b11111000100111000;
mem[353]=17'b00000000001101010;
mem[354]=17'b11111111111101011;
mem[355]=17'b11101111110101011;
mem[356]=17'b11111111111011011;
mem[357]=17'b11111111111110100;
mem[358]=17'b11110010001111101;
mem[359]=17'b00000010011110111;
mem[360]=17'b11111111000011101;
mem[361]=17'b00000111101000001;
mem[362]=17'b11111111011100000;
mem[363]=17'b00000001101000000;
mem[364]=17'b00000001001100110;
mem[365]=17'b00000011110100111;
mem[366]=17'b00000011010010100;
mem[367]=17'b11111000100001111;
mem[368]=17'b11111100000011100;
mem[369]=17'b00000001010101101;
mem[370]=17'b00000000001001100;
mem[371]=17'b00000000001111000;
mem[372]=17'b00000110111111110;
mem[373]=17'b00000000000111010;
mem[374]=17'b11111101101110111;
mem[375]=17'b11111110101011010;
mem[376]=17'b11111110011001100;
mem[377]=17'b00000000010010001;
mem[378]=17'b11111111011100100;
mem[379]=17'b11111111101101001;
mem[380]=17'b11111011001111000;
mem[381]=17'b00000001011000110;
mem[382]=17'b00000001101001111;
mem[383]=17'b11111101111010011;
mem[384]=17'b00000001011100001;
mem[385]=17'b11111111011011100;
mem[386]=17'b00000000001000110;
mem[387]=17'b00000001100101110;
mem[388]=17'b11111111110000100;
mem[389]=17'b00000001100101101;
mem[390]=17'b00000000011111100;
mem[391]=17'b11111110110010110;
mem[392]=17'b11111111101111011;
mem[393]=17'b00000000000010110;
mem[394]=17'b00000000010010110;
mem[395]=17'b11111111110101101;
mem[396]=17'b11111111101110011;
mem[397]=17'b11111010011010100;
mem[398]=17'b11111111111010000;
mem[399]=17'b11111111000000010;
mem[400]=17'b00000000011000000;
mem[401]=17'b11111100001100000;
mem[402]=17'b11111111000100000;
mem[403]=17'b00000001001100100;
mem[404]=17'b11111001010101110;
mem[405]=17'b00010010001001100;
mem[406]=17'b00000000001011111;
mem[407]=17'b00000010111110101;
mem[408]=17'b00000000000111111;
mem[409]=17'b11110101110111100;
mem[410]=17'b00000000001000110;
mem[411]=17'b00000001101011001;
mem[412]=17'b11111111101111100;
mem[413]=17'b11110111100111010;
mem[414]=17'b11111011010010111;
mem[415]=17'b00001000001010111;
mem[416]=17'b11111010111010111;
mem[417]=17'b11111111111010110;
mem[418]=17'b00000100010111010;
mem[419]=17'b00000010110100101;
mem[420]=17'b00000000000000110;
mem[421]=17'b11111110011010011;
mem[422]=17'b11111110100011110;
mem[423]=17'b00000000100001000;
mem[424]=17'b00011010110100011;
mem[425]=17'b00000000011101011;
mem[426]=17'b11111111100100100;
mem[427]=17'b11111111000001001;
mem[428]=17'b00000000010100110;
mem[429]=17'b00000000000100010;
mem[430]=17'b11111010101010011;
mem[431]=17'b11111001111000111;
mem[432]=17'b00000000100100011;
mem[433]=17'b11111000110000100;
mem[434]=17'b11111111100001010;
mem[435]=17'b11111111110110001;
mem[436]=17'b00000000000011110;
mem[437]=17'b11111110110000010;
mem[438]=17'b11111010101111110;
mem[439]=17'b00000001000100000;
mem[440]=17'b11111111001011011;
mem[441]=17'b00000000101001100;
mem[442]=17'b11111100101110101;
mem[443]=17'b00000000000100000;
mem[444]=17'b00000000001000001;
mem[445]=17'b11111110011011000;
mem[446]=17'b00001001101010101;
mem[447]=17'b11111111110110100;
mem[448]=17'b11111111100000001;
mem[449]=17'b11111111100011011;
mem[450]=17'b11111111101001000;
mem[451]=17'b00000001110000011;
mem[452]=17'b00000000101110111;
mem[453]=17'b11111000111011110;
mem[454]=17'b11111111110111010;
mem[455]=17'b11111111010100101;
mem[456]=17'b00000000001100100;
mem[457]=17'b11110101111110000;
mem[458]=17'b11111111100011011;
mem[459]=17'b00000000001001100;
mem[460]=17'b11111111110100001;
mem[461]=17'b00000011011111111;
mem[462]=17'b11111111101100101;
mem[463]=17'b00000000001001111;
mem[464]=17'b11111110000000001;
mem[465]=17'b11111111110001111;
mem[466]=17'b00000000001101010;
mem[467]=17'b00000000001000101;
mem[468]=17'b11111111110111011;
mem[469]=17'b00000000000011010;
mem[470]=17'b00000000000110100;
mem[471]=17'b00000000001010111;
mem[472]=17'b11111111101000010;
mem[473]=17'b11111111101100111;
mem[474]=17'b00000000011110000;
mem[475]=17'b11111111111100011;
mem[476]=17'b00000001110010011;
mem[477]=17'b11111100001000101;
mem[478]=17'b11111111111101100;
mem[479]=17'b00000000011011000;
mem[480]=17'b11111111101001011;
mem[481]=17'b00000000110110000;
mem[482]=17'b11111101001000000;
mem[483]=17'b11111100111011101;
mem[484]=17'b00000000000000001;
mem[485]=17'b11111110001011010;
mem[486]=17'b00000000011100110;
mem[487]=17'b11111111000000100;
mem[488]=17'b11111101011011111;
mem[489]=17'b11111110001000001;
mem[490]=17'b00000000101001100;
mem[491]=17'b11111101101010000;
mem[492]=17'b00000000000000010;
mem[493]=17'b11111111111111110;
mem[494]=17'b00000001000001001;
mem[495]=17'b00000101011111000;
mem[496]=17'b11111110101110000;
mem[497]=17'b00000000101010110;
mem[498]=17'b11101111011110011;
mem[499]=17'b00000000001101001;
mem[500]=17'b11111111101011010;
mem[501]=17'b00000000011111011;
mem[502]=17'b11111111110011011;
mem[503]=17'b00000011000101001;
mem[504]=17'b00000000001111000;
mem[505]=17'b11111010011101100;
mem[506]=17'b11111010000110011;
mem[507]=17'b00000000000101110;
mem[508]=17'b00000001011011110;
mem[509]=17'b11110001001010100;
mem[510]=17'b11111100100011010;
mem[511]=17'b00000010111110000;
mem[512]=17'b00000010000000000;
mem[513]=17'b00000000011001110;
mem[514]=17'b00000000010011010;
mem[515]=17'b00000000101000001;
mem[516]=17'b11111110111110010;
mem[517]=17'b11111111000110110;
mem[518]=17'b00000000011001000;
mem[519]=17'b00000001000101011;
mem[520]=17'b00000000000110010;
mem[521]=17'b00000001110111111;
mem[522]=17'b00000000000111101;
mem[523]=17'b00000000000111010;
mem[524]=17'b00000100111011011;
mem[525]=17'b11111101111100011;
mem[526]=17'b00000000011010011;
mem[527]=17'b11111110111111011;
mem[528]=17'b11111110110110010;
mem[529]=17'b11111111111010010;
mem[530]=17'b11111111110110011;
mem[531]=17'b11111111101001011;
mem[532]=17'b11111110010010100;
mem[533]=17'b00000000010110000;
mem[534]=17'b11111010010111001;
mem[535]=17'b11111111101001010;
mem[536]=17'b00000000000100001;
mem[537]=17'b00000000100001110;
mem[538]=17'b11111111100101000;
mem[539]=17'b11111101000011000;
mem[540]=17'b11111100101000111;
mem[541]=17'b11111110101111000;
mem[542]=17'b11111111111111100;
mem[543]=17'b11111111110011000;
mem[544]=17'b11111111100010011;
mem[545]=17'b01101010011011110;
mem[546]=17'b11011110101101110;
mem[547]=17'b00010110100000011;
mem[548]=17'b00000001110111000;
mem[549]=17'b11111111000100111;
mem[550]=17'b11101001110001001;
mem[551]=17'b11111101110100110;
mem[552]=17'b00000001001010111;
mem[553]=17'b00001010111110001;
mem[554]=17'b11111101110000110;
mem[555]=17'b00000000111000011;
mem[556]=17'b11110011010001001;
mem[557]=17'b11111110000010100;
mem[558]=17'b11111111100100010;
mem[559]=17'b11111101010101101;
mem[560]=17'b00000000100000100;
mem[561]=17'b00000010011010000;
mem[562]=17'b11111011110111001;
mem[563]=17'b00000101100001011;
mem[564]=17'b00000000001111110;
mem[565]=17'b11111000011101111;
mem[566]=17'b11111111101001000;
mem[567]=17'b00000000111000101;
mem[568]=17'b11111111100001101;
mem[569]=17'b00000000011101010;
mem[570]=17'b00000000001100101;
mem[571]=17'b00000000001001111;
mem[572]=17'b11111111110001100;
mem[573]=17'b11111111111110000;
mem[574]=17'b00000000000000011;
mem[575]=17'b00000001101101110;
mem[576]=17'b11111111111100110;
mem[577]=17'b11111110110001100;
mem[578]=17'b11111011011000100;
mem[579]=17'b11111101001001110;
mem[580]=17'b00000011111001011;
mem[581]=17'b11111111110011101;
mem[582]=17'b00000000101000010;
mem[583]=17'b11111111111101110;
mem[584]=17'b11111110110010111;
mem[585]=17'b00000000000101101;
mem[586]=17'b00000000011100111;
mem[587]=17'b00001010001110100;
mem[588]=17'b11111100011100011;
mem[589]=17'b11111111000000100;
mem[590]=17'b00000000011010011;
mem[591]=17'b00000001011111001;
mem[592]=17'b11111111010001101;
mem[593]=17'b11111110111011100;
mem[594]=17'b00011101000011111;
mem[595]=17'b00000000011111001;
mem[596]=17'b11111111011000000;
mem[597]=17'b00000000010110111;
mem[598]=17'b00000111010000000;
mem[599]=17'b11111110111101111;
mem[600]=17'b00000000001000010;
mem[601]=17'b11111010101101001;
mem[602]=17'b11111111011001001;
mem[603]=17'b00000000101111010;
mem[604]=17'b11111111111011011;
mem[605]=17'b11110111101110011;
mem[606]=17'b11111111110010101;
mem[607]=17'b11111111100100011;
mem[608]=17'b11111111111000110;
mem[609]=17'b00100010110000000;
mem[610]=17'b11111111011010111;
mem[611]=17'b00000000001111101;
mem[612]=17'b11111111111001001;
mem[613]=17'b11111110010101100;
mem[614]=17'b11111111111110110;
mem[615]=17'b00000110001111011;
mem[616]=17'b00000001100101000;
mem[617]=17'b11111111001000010;
mem[618]=17'b00000001100010010;
mem[619]=17'b11111010111010100;
mem[620]=17'b00000000001010011;
mem[621]=17'b00000000100101011;
mem[622]=17'b00000000000000100;
mem[623]=17'b00000000010000110;
mem[624]=17'b00000000010100010;
mem[625]=17'b11111011101100011;
mem[626]=17'b00000010110111011;
mem[627]=17'b11111110010100110;
mem[628]=17'b00000001110101101;
mem[629]=17'b11111110110101010;
mem[630]=17'b11110101000011110;
mem[631]=17'b00000001110100101;
mem[632]=17'b11111100111000110;
mem[633]=17'b11111111111110100;
mem[634]=17'b00000000001111101;
mem[635]=17'b11111111110000100;
mem[636]=17'b11111111010101100;
mem[637]=17'b11111101010110000;
mem[638]=17'b11111111010100110;
mem[639]=17'b11010100000101111;
mem[640]=17'b00000000111110110;
mem[641]=17'b11111111111101101;
mem[642]=17'b11111110111101010;
mem[643]=17'b11111111110001111;
mem[644]=17'b00000000111000010;
mem[645]=17'b00011000100110010;
mem[646]=17'b11111101100010100;
mem[647]=17'b00000000110101000;
mem[648]=17'b11111111010010101;
mem[649]=17'b11111100001010000;
mem[650]=17'b00000000010010011;
mem[651]=17'b11111110101001011;
mem[652]=17'b00000001011001110;
mem[653]=17'b00000001000101001;
mem[654]=17'b00000000001011100;
mem[655]=17'b00000010010010110;
mem[656]=17'b11111110101010010;
mem[657]=17'b11111111100101111;
mem[658]=17'b11111110000000001;
mem[659]=17'b11111000110111001;
mem[660]=17'b00000000000101110;
mem[661]=17'b11110101001001100;
mem[662]=17'b00000001001101100;
mem[663]=17'b11111110101101001;
mem[664]=17'b11111111101101000;
mem[665]=17'b00000000000000001;
mem[666]=17'b11111110100011100;
mem[667]=17'b11111111001100000;
mem[668]=17'b00000110000101111;
mem[669]=17'b11111110011001000;
mem[670]=17'b00000111111001101;
mem[671]=17'b00000001101100001;
mem[672]=17'b11111111110001001;
mem[673]=17'b00000000100011111;
mem[674]=17'b00000000000110000;
mem[675]=17'b00000010010110010;
mem[676]=17'b00000000101000101;
mem[677]=17'b00000000001000111;
mem[678]=17'b00000011011010010;
mem[679]=17'b00000100010111100;
mem[680]=17'b00000000000011001;
mem[681]=17'b00000001101010100;
mem[682]=17'b00000000000111010;
mem[683]=17'b00000000001000100;
mem[684]=17'b00000000000000011;
mem[685]=17'b11111110110101001;
mem[686]=17'b00000001101100111;
mem[687]=17'b11110010000010011;
mem[688]=17'b11111111110101000;
mem[689]=17'b00000000001100011;
mem[690]=17'b11111111111111111;
mem[691]=17'b00001001101011110;
mem[692]=17'b00000000010000111;
mem[693]=17'b00000000000000001;
mem[694]=17'b11111111011101010;
mem[695]=17'b00000000100101011;
mem[696]=17'b11111111100110110;
mem[697]=17'b11111111001100111;
mem[698]=17'b11111111001000011;
mem[699]=17'b00000000010001010;
mem[700]=17'b00000011101110000;
mem[701]=17'b11111111101000010;
mem[702]=17'b00000000011101010;
mem[703]=17'b00000000000011110;
mem[704]=17'b00000000101101011;
mem[705]=17'b00000001111011000;
mem[706]=17'b11111110101111110;
mem[707]=17'b00000000101100010;
mem[708]=17'b11111111101111010;
mem[709]=17'b00000000100010011;
mem[710]=17'b00000000110010000;
mem[711]=17'b11111101001010010;
mem[712]=17'b00000000001001001;
mem[713]=17'b00000000010101010;
mem[714]=17'b00000000101011000;
mem[715]=17'b00000010100011110;
mem[716]=17'b00000000101011011;
mem[717]=17'b00000000111100010;
mem[718]=17'b00000000010010111;
mem[719]=17'b11111110100110100;
mem[720]=17'b00000011001100000;
mem[721]=17'b00000001100001110;
mem[722]=17'b00000001010110001;
mem[723]=17'b11111101011011100;
mem[724]=17'b11111111111000001;
mem[725]=17'b11111111111001011;
mem[726]=17'b00000010001101110;
mem[727]=17'b11111000101010000;
mem[728]=17'b11111111111100100;
mem[729]=17'b11111111011100111;
mem[730]=17'b00000010000000100;
mem[731]=17'b11111110010111110;
mem[732]=17'b11111110101000000;
mem[733]=17'b11111111111111111;
mem[734]=17'b00000000010011110;
mem[735]=17'b11111110101001010;
mem[736]=17'b00000000000010110;
mem[737]=17'b00000000000011111;
mem[738]=17'b00000001000101110;
mem[739]=17'b11111111111100110;
mem[740]=17'b11111100100000110;
mem[741]=17'b11110110111011101;
mem[742]=17'b00000000011000100;
mem[743]=17'b11111110110011000;
mem[744]=17'b11111111001100000;
mem[745]=17'b00000000000101000;
mem[746]=17'b11111110101100011;
mem[747]=17'b00000000101100100;
mem[748]=17'b11111101010000110;
mem[749]=17'b11111100100010000;
mem[750]=17'b11111111001011110;
mem[751]=17'b11111110000110111;
mem[752]=17'b00000000010101110;
mem[753]=17'b00000001111001010;
mem[754]=17'b11111111000011011;
mem[755]=17'b00000001010100001;
mem[756]=17'b11111111100100010;
mem[757]=17'b00000010111011101;
mem[758]=17'b00000000000010001;
mem[759]=17'b11111011101001000;
mem[760]=17'b11101101000011100;
mem[761]=17'b00000001000111011;
mem[762]=17'b00000000011000111;
mem[763]=17'b00000010011011100;
mem[764]=17'b11111110011111111;
mem[765]=17'b11110001101010110;
mem[766]=17'b11101110010101111;
mem[767]=17'b00000110001101100;
mem[768]=17'b00001001010100110;
mem[769]=17'b11111101100100000;
mem[770]=17'b00000010100110100;
mem[771]=17'b11111111010011011;
mem[772]=17'b11111111111111100;
mem[773]=17'b11101010000100011;
mem[774]=17'b11111111110100100;
mem[775]=17'b00000000001001000;
mem[776]=17'b11111111011000000;
mem[777]=17'b00000000011110111;
mem[778]=17'b00000000000101101;
mem[779]=17'b11111111111101001;
mem[780]=17'b11110110100111110;
mem[781]=17'b11111111101101011;
mem[782]=17'b00000001000111001;
mem[783]=17'b00000000001001010;
mem[784]=17'b00000000010001000;
mem[785]=17'b00000000000011000;
mem[786]=17'b11111111011001000;
mem[787]=17'b11111111110111010;
mem[788]=17'b00000000010010110;
mem[789]=17'b00000000000100000;
mem[790]=17'b00000000001001011;
mem[791]=17'b00000000110001000;
mem[792]=17'b11111100111010010;
mem[793]=17'b00000000100010010;
mem[794]=17'b00000000100100001;
mem[795]=17'b11111111001101101;
mem[796]=17'b00000000100010110;
mem[797]=17'b00000001001011100;
mem[798]=17'b11111111001010000;
mem[799]=17'b00000000110100001;
mem[800]=17'b00000010000001111;
mem[801]=17'b11111111111101101;
mem[802]=17'b11111111000001100;
mem[803]=17'b00000101001110110;
mem[804]=17'b00000000000110001;
mem[805]=17'b00000010010000001;
mem[806]=17'b11111111011100001;
mem[807]=17'b11111110111000010;
mem[808]=17'b00000001101101101;
mem[809]=17'b11111111111011001;
mem[810]=17'b11111111111101110;
mem[811]=17'b00000001010011010;
mem[812]=17'b11111111111111010;
mem[813]=17'b00000001011001100;
mem[814]=17'b11111111000100010;
mem[815]=17'b00000010010100010;
mem[816]=17'b00000010100110100;
mem[817]=17'b11111111110010000;
mem[818]=17'b00000000000111101;
mem[819]=17'b11111101000110100;
mem[820]=17'b11111110111100001;
mem[821]=17'b11111111110101101;
mem[822]=17'b11111100001011111;
mem[823]=17'b00000000000100100;
mem[824]=17'b00000000011001001;
mem[825]=17'b00000001011000100;
mem[826]=17'b00000000100110001;
mem[827]=17'b11111110110000011;
mem[828]=17'b00000010101010111;
mem[829]=17'b00000110101100110;
mem[830]=17'b11111111011111101;
mem[831]=17'b11111111101111101;
mem[832]=17'b00000001011010011;
mem[833]=17'b00000000001100011;
mem[834]=17'b00000000110010101;
mem[835]=17'b11111011100101110;
mem[836]=17'b11111111110111100;
mem[837]=17'b11111111110111100;
mem[838]=17'b00000000001001100;
mem[839]=17'b00000000011100011;
mem[840]=17'b11111110111010110;
mem[841]=17'b11111111111111111;
mem[842]=17'b00000000000010111;
mem[843]=17'b00000000110110111;
mem[844]=17'b00000001001011101;
mem[845]=17'b00000010100101001;
mem[846]=17'b00000000111100001;
mem[847]=17'b00000010000101101;
mem[848]=17'b00000000100110111;
mem[849]=17'b11111111111000001;
mem[850]=17'b11111111010100010;
mem[851]=17'b11111110001000011;
mem[852]=17'b00001010011101111;
mem[853]=17'b00000000101101110;
mem[854]=17'b00000000001001001;
mem[855]=17'b11111101111001100;
mem[856]=17'b00000001100011000;
mem[857]=17'b11111111001000110;
mem[858]=17'b11111111011111011;
mem[859]=17'b00000000000001010;
mem[860]=17'b00000000000000000;
mem[861]=17'b11111111101010101;
mem[862]=17'b00000000111111000;
mem[863]=17'b00000000111000001;
mem[864]=17'b11111100011100010;
mem[865]=17'b00000000011010001;
mem[866]=17'b00000101111110100;
mem[867]=17'b00000000010011110;
mem[868]=17'b00000000010011001;
mem[869]=17'b00000000001100010;
mem[870]=17'b00000000000110010;
mem[871]=17'b11111111011101001;
mem[872]=17'b00000000011101011;
mem[873]=17'b00110010010011011;
mem[874]=17'b11111111000100110;
mem[875]=17'b11110111111010100;
mem[876]=17'b00000000000000001;
mem[877]=17'b11111111111101000;
mem[878]=17'b00000100101110110;
mem[879]=17'b11111110010111110;
mem[880]=17'b11111111010000110;
mem[881]=17'b11111110101001011;
mem[882]=17'b00000000110110100;
mem[883]=17'b00000000010110110;
mem[884]=17'b00000000010101011;
mem[885]=17'b00000000001111000;
mem[886]=17'b00000000001011001;
mem[887]=17'b00000000001001110;
mem[888]=17'b00000000000010000;
mem[889]=17'b11111011101100110;
mem[890]=17'b00000000000001101;
mem[891]=17'b00000100011001011;
mem[892]=17'b11111111110101110;
mem[893]=17'b11111110010110001;
mem[894]=17'b00000000101111001;
mem[895]=17'b11111110011010010;
mem[896]=17'b00000000010011101;
mem[897]=17'b11111101001100010;
mem[898]=17'b00000000010010010;
mem[899]=17'b11111001001100101;
mem[900]=17'b11111101100110001;
mem[901]=17'b00011010101000100;
mem[902]=17'b11111111101100101;
mem[903]=17'b11111111110100000;
mem[904]=17'b00000101100010110;
mem[905]=17'b00000000100111101;
mem[906]=17'b00001111100100100;
mem[907]=17'b11111100110101001;
mem[908]=17'b11111111000000011;
mem[909]=17'b11111111110011100;
mem[910]=17'b11111111100000100;
mem[911]=17'b11111110101001001;
mem[912]=17'b00000110100001011;
mem[913]=17'b11111111111000101;
mem[914]=17'b11111010000100110;
mem[915]=17'b00001001010011110;
mem[916]=17'b00000001100101110;
mem[917]=17'b00000000001000101;
mem[918]=17'b11111111111101101;
mem[919]=17'b11111111111100101;
mem[920]=17'b00000000100011100;
mem[921]=17'b11111111111010001;
mem[922]=17'b11111111111111101;
mem[923]=17'b00000000001001111;
mem[924]=17'b11111111001001101;
mem[925]=17'b11111111111100111;
mem[926]=17'b11111111111110001;
mem[927]=17'b00000000001111001;
mem[928]=17'b00000000011110101;
mem[929]=17'b11111111101100011;
mem[930]=17'b11111110100100000;
mem[931]=17'b11111111111010110;
mem[932]=17'b00000000111000110;
mem[933]=17'b00000000100010000;
mem[934]=17'b11111111101100100;
mem[935]=17'b11111111000011011;
mem[936]=17'b11111101000010010;
mem[937]=17'b00000000001011110;
mem[938]=17'b00010000101101001;
mem[939]=17'b11111111110110011;
mem[940]=17'b00000001111101111;
mem[941]=17'b11111111101011101;
mem[942]=17'b00000000000000011;
mem[943]=17'b00000101111110001;
mem[944]=17'b00000010010000111;
mem[945]=17'b11111110001111101;
mem[946]=17'b00000000110111110;
mem[947]=17'b00000000110101100;
mem[948]=17'b11111111111010010;
mem[949]=17'b11111111010000100;
mem[950]=17'b11111010111100001;
mem[951]=17'b11111111111011101;
mem[952]=17'b11111111110101011;
mem[953]=17'b00000011011101001;
mem[954]=17'b11111110101110101;
mem[955]=17'b00000000001101001;
mem[956]=17'b00000000001100111;
mem[957]=17'b11111101111100001;
mem[958]=17'b00000001000101111;
mem[959]=17'b11111111110100011;
mem[960]=17'b00000000011110100;
mem[961]=17'b11111110011111011;
mem[962]=17'b11111111110110010;
mem[963]=17'b11111110010000100;
mem[964]=17'b11111101111100001;
mem[965]=17'b11111111100101010;
mem[966]=17'b00000001010111001;
mem[967]=17'b11111111110010010;
mem[968]=17'b00000000011011100;
mem[969]=17'b00000110010110010;
mem[970]=17'b11110000010100110;
mem[971]=17'b00000001001001011;
mem[972]=17'b11111111011010111;
mem[973]=17'b11111111011110010;
mem[974]=17'b11101010000110100;
mem[975]=17'b00000000000000111;
mem[976]=17'b11111111111001101;
mem[977]=17'b11111111110101100;
mem[978]=17'b11111111111111010;
mem[979]=17'b00000001010111000;
mem[980]=17'b00000000010110000;
mem[981]=17'b11111111111110011;
mem[982]=17'b11111111000010101;
mem[983]=17'b11111111011111100;
mem[984]=17'b11111111101101110;
mem[985]=17'b11111010111110010;
mem[986]=17'b11111111001110010;
mem[987]=17'b00000000111000010;
mem[988]=17'b00000100111011111;
mem[989]=17'b00000111100111000;
mem[990]=17'b00000001100101101;
mem[991]=17'b11111111101100110;
mem[992]=17'b00000001010010001;
mem[993]=17'b11111111011001111;
mem[994]=17'b11111111110110100;
mem[995]=17'b11111101111010000;
mem[996]=17'b00000001110111100;
mem[997]=17'b00000101100101100;
mem[998]=17'b00000001011111000;
mem[999]=17'b11111011010010001;
mem[1000]=17'b00000000001110101;
mem[1001]=17'b11111111111010100;
mem[1002]=17'b00000010001000010;
mem[1003]=17'b11111111111011000;
mem[1004]=17'b11111111111110011;
mem[1005]=17'b11111111100110010;
mem[1006]=17'b00000000011111110;
mem[1007]=17'b00000000010111010;
mem[1008]=17'b11111100101010111;
mem[1009]=17'b00000000001010010;
mem[1010]=17'b00000000101011101;
mem[1011]=17'b11111111111011011;
mem[1012]=17'b11101000101111011;
mem[1013]=17'b11111101000100000;
mem[1014]=17'b00000000011100000;
mem[1015]=17'b11111111111010000;
mem[1016]=17'b00000001010011011;
mem[1017]=17'b00000100010000101;
mem[1018]=17'b00000000101000110;
mem[1019]=17'b00000000001011100;
mem[1020]=17'b11111110111101110;
mem[1021]=17'b11111111001000000;
mem[1022]=17'b00000000100001101;
mem[1023]=17'b11111111100101111;
mem[1024]=17'b00001101111001011;
mem[1025]=17'b00000100110011110;
mem[1026]=17'b00000000100111110;
mem[1027]=17'b11111111110000000;
mem[1028]=17'b11111111110010111;
mem[1029]=17'b11111110001110010;
mem[1030]=17'b11111111111000010;
mem[1031]=17'b11111110110110010;
mem[1032]=17'b00000000010111101;
mem[1033]=17'b11101100000010101;
mem[1034]=17'b10111001101111101;
mem[1035]=17'b11110110111100111;
mem[1036]=17'b00001110010010111;
mem[1037]=17'b00000000011100000;
mem[1038]=17'b11111111111000100;
mem[1039]=17'b00000000010101011;
mem[1040]=17'b11111111100011110;
mem[1041]=17'b00000000000001011;
mem[1042]=17'b11111110100011111;
mem[1043]=17'b00000000001011011;
mem[1044]=17'b00000000000010100;
mem[1045]=17'b00000000000110101;
mem[1046]=17'b00000000001100000;
mem[1047]=17'b00000000000001001;
mem[1048]=17'b00000000011011111;
mem[1049]=17'b11111111110101000;
mem[1050]=17'b11111101010110101;
mem[1051]=17'b00000000000101100;
mem[1052]=17'b11111011000010000;
mem[1053]=17'b00000001001110100;
mem[1054]=17'b00000001010010100;
mem[1055]=17'b00000000001000001;
mem[1056]=17'b00000000010001111;
mem[1057]=17'b00000000000011110;
mem[1058]=17'b00000000000001010;
mem[1059]=17'b11111110111111000;
mem[1060]=17'b11111100000110000;
mem[1061]=17'b00000000000000000;
mem[1062]=17'b11111111010001111;
mem[1063]=17'b00000000011010011;
mem[1064]=17'b11111111111010001;
mem[1065]=17'b00000000001001101;
mem[1066]=17'b11111111110011100;
mem[1067]=17'b11111100000000111;
mem[1068]=17'b00000000110000001;
mem[1069]=17'b11111110000111001;
mem[1070]=17'b00000000100101110;
mem[1071]=17'b00000001110100100;
mem[1072]=17'b00000000010111010;
mem[1073]=17'b00000010111100000;
mem[1074]=17'b11111101000111111;
mem[1075]=17'b11111100001101000;
mem[1076]=17'b00000000001110110;
mem[1077]=17'b00000010001011111;
mem[1078]=17'b11111101000000111;
mem[1079]=17'b11111111111100010;
mem[1080]=17'b00000000110101010;
mem[1081]=17'b11111110101110010;
mem[1082]=17'b00000000111001101;
mem[1083]=17'b11111110001010010;
mem[1084]=17'b00010000010000111;
mem[1085]=17'b11100001110101111;
mem[1086]=17'b00000000101010011;
mem[1087]=17'b00000000001001111;
mem[1088]=17'b00000000001000101;
mem[1089]=17'b00000001000100101;
mem[1090]=17'b00000000000001001;
mem[1091]=17'b11100110111011110;
mem[1092]=17'b11111110111100111;
mem[1093]=17'b11111110011011110;
mem[1094]=17'b11111111110001101;
mem[1095]=17'b00000000010110100;
mem[1096]=17'b11111111110101101;
mem[1097]=17'b11111111001110100;
mem[1098]=17'b00000000010011011;
mem[1099]=17'b01101101001011000;
mem[1100]=17'b00000011001000010;
mem[1101]=17'b11111101101001111;
mem[1102]=17'b11111110110001000;
mem[1103]=17'b00000000011100101;
mem[1104]=17'b11111110111101101;
mem[1105]=17'b11111011001111001;
mem[1106]=17'b00000000001101001;
mem[1107]=17'b11111101111111000;
mem[1108]=17'b00000000100001011;
mem[1109]=17'b00000000000110111;
mem[1110]=17'b00000001000100011;
mem[1111]=17'b11111111101100100;
mem[1112]=17'b11101111111000001;
mem[1113]=17'b00000100011100000;
mem[1114]=17'b00000001011101100;
mem[1115]=17'b11111110101110000;
mem[1116]=17'b11111111110110010;
mem[1117]=17'b00000000001001110;
mem[1118]=17'b00000000000111110;
mem[1119]=17'b11111110111111111;
mem[1120]=17'b11111110010000111;
mem[1121]=17'b11111100101110010;
mem[1122]=17'b00000000000101001;
mem[1123]=17'b11111111011111110;
mem[1124]=17'b00000000000110100;
mem[1125]=17'b00000000011001001;
mem[1126]=17'b00000000000111001;
mem[1127]=17'b11111111110111011;
mem[1128]=17'b00000001011101010;
mem[1129]=17'b11111100100000101;
mem[1130]=17'b11111010111010101;
mem[1131]=17'b11111111101100000;
mem[1132]=17'b00000010010010011;
mem[1133]=17'b11111111110111100;
mem[1134]=17'b00000001110111010;
mem[1135]=17'b00000000000001101;
mem[1136]=17'b11111110011011001;
mem[1137]=17'b11111110110101111;
mem[1138]=17'b11111111111011001;
mem[1139]=17'b11111111100111011;
mem[1140]=17'b00000001101011110;
mem[1141]=17'b00000001101000100;
mem[1142]=17'b00000000000110001;
mem[1143]=17'b11111111011101010;
mem[1144]=17'b11111101100000000;
mem[1145]=17'b11111011001001010;
mem[1146]=17'b11111111011010001;
mem[1147]=17'b11111101011111110;
mem[1148]=17'b11111111110011001;
mem[1149]=17'b11111111100100110;
mem[1150]=17'b00000011111010011;
mem[1151]=17'b11101100100100101;
mem[1152]=17'b00000000111001100;
mem[1153]=17'b00000001010001100;
mem[1154]=17'b11111110001100000;
mem[1155]=17'b11111110111011100;
mem[1156]=17'b11111101110100001;
mem[1157]=17'b00000001101001011;
mem[1158]=17'b11111111110011010;
mem[1159]=17'b00000000110100010;
mem[1160]=17'b00011110111110001;
mem[1161]=17'b00000000000010101;
mem[1162]=17'b00000000000100010;
mem[1163]=17'b11111101110101101;
mem[1164]=17'b00001001001000011;
mem[1165]=17'b00000000010000000;
mem[1166]=17'b11100111111110001;
mem[1167]=17'b11111111111110110;
mem[1168]=17'b11010110100110000;
mem[1169]=17'b00000000000001101;
mem[1170]=17'b00000000000100111;
mem[1171]=17'b11111111011010101;
mem[1172]=17'b00000000001010101;
mem[1173]=17'b11111111100111101;
mem[1174]=17'b00000001110010100;
mem[1175]=17'b00000010100111011;
mem[1176]=17'b11010101101011101;
mem[1177]=17'b00000000101000010;
mem[1178]=17'b00000000000101000;
mem[1179]=17'b11111111101110011;
mem[1180]=17'b11111111111000101;
mem[1181]=17'b11111111100001100;
mem[1182]=17'b00000101011101000;
mem[1183]=17'b11111111001111111;
mem[1184]=17'b11111111101101000;
mem[1185]=17'b11111100100001000;
mem[1186]=17'b11111100111100100;
mem[1187]=17'b00000110011001100;
mem[1188]=17'b11111111001111001;
mem[1189]=17'b11111110010011000;
mem[1190]=17'b00000000001011100;
mem[1191]=17'b00000010000100011;
mem[1192]=17'b00000001100101000;
mem[1193]=17'b00000000010100101;
mem[1194]=17'b11111111111001000;
mem[1195]=17'b00000000010011101;
mem[1196]=17'b11111111110010111;
mem[1197]=17'b00000000001001111;
mem[1198]=17'b00011100101000111;
mem[1199]=17'b11111110100001100;
mem[1200]=17'b11111111111000000;
mem[1201]=17'b00000000001010000;
mem[1202]=17'b11111101100011100;
mem[1203]=17'b00000000101101010;
mem[1204]=17'b11111111110010100;
mem[1205]=17'b00000000000000001;
mem[1206]=17'b00000001000011001;
mem[1207]=17'b11111110010110101;
mem[1208]=17'b00000000000000010;
mem[1209]=17'b11111111001111010;
mem[1210]=17'b00000000001110001;
mem[1211]=17'b11111110110110010;
mem[1212]=17'b11111111011001100;
mem[1213]=17'b11111111110101001;
mem[1214]=17'b00000010001101011;
mem[1215]=17'b00001000100001010;
mem[1216]=17'b11111111011000101;
mem[1217]=17'b11111110111001111;
mem[1218]=17'b00000000101000110;
mem[1219]=17'b00000000000100100;
mem[1220]=17'b11111111001100000;
mem[1221]=17'b11111101000101010;
mem[1222]=17'b11111111111110100;
mem[1223]=17'b11111111110111001;
mem[1224]=17'b00000000000000001;
mem[1225]=17'b00000001110011100;
mem[1226]=17'b11111110011000111;
mem[1227]=17'b00000101001101100;
mem[1228]=17'b00000011011101101;
mem[1229]=17'b00000100100010001;
mem[1230]=17'b11111111100100000;
mem[1231]=17'b11111110000110001;
mem[1232]=17'b00000001100111100;
mem[1233]=17'b11110001011011010;
mem[1234]=17'b11111110100111110;
mem[1235]=17'b11111101101111011;
mem[1236]=17'b00001011111011000;
mem[1237]=17'b11111111011011011;
mem[1238]=17'b00000000111001010;
mem[1239]=17'b11111111101001101;
mem[1240]=17'b00001000000010000;
mem[1241]=17'b00000000000100011;
mem[1242]=17'b00000000100001111;
mem[1243]=17'b11111110001111110;
mem[1244]=17'b11111110111001100;
mem[1245]=17'b00000000001000110;
mem[1246]=17'b00000000000111001;
mem[1247]=17'b00000000011110111;
mem[1248]=17'b11111111101100000;
mem[1249]=17'b11111111010000111;
mem[1250]=17'b11111111111100010;
mem[1251]=17'b00000000000101011;
mem[1252]=17'b11111111000001101;
mem[1253]=17'b00000000000011011;
mem[1254]=17'b00000000000010101;
mem[1255]=17'b00001001101100110;
mem[1256]=17'b11111111000110010;
mem[1257]=17'b11111101100010110;
mem[1258]=17'b00000000000110001;
mem[1259]=17'b00000110000111000;
mem[1260]=17'b11111111111110001;
mem[1261]=17'b00000000011111111;
mem[1262]=17'b11111101100001101;
mem[1263]=17'b11111110111110011;
mem[1264]=17'b00000000000110101;
mem[1265]=17'b00011110000111101;
mem[1266]=17'b00000001100010101;
mem[1267]=17'b00000001111000111;
mem[1268]=17'b00000000000011001;
mem[1269]=17'b11111111010101110;
mem[1270]=17'b00000000001001011;
mem[1271]=17'b00001000110100011;
mem[1272]=17'b00000000101011000;
mem[1273]=17'b11111111001101001;
mem[1274]=17'b00000000100011011;
mem[1275]=17'b11111111111101000;
mem[1276]=17'b00000000000110010;
mem[1277]=17'b11111111111011001;
mem[1278]=17'b11110101111111011;
mem[1279]=17'b11111000101011001;
mem[1280]=17'b00000000011111000;
mem[1281]=17'b00000000011001000;
mem[1282]=17'b11111111101001101;
mem[1283]=17'b00000010110010101;
mem[1284]=17'b11111111111101010;
mem[1285]=17'b11111111101100110;
mem[1286]=17'b11111111001000010;
mem[1287]=17'b00001101000010000;
mem[1288]=17'b11111111100001111;
mem[1289]=17'b00000011000001111;
mem[1290]=17'b11111011011011101;
mem[1291]=17'b00000000111110100;
mem[1292]=17'b00000000010110100;
mem[1293]=17'b11111111101111100;
mem[1294]=17'b00000010001011111;
mem[1295]=17'b00000000000000011;
mem[1296]=17'b11111110101011110;
mem[1297]=17'b00000000101001101;
mem[1298]=17'b11111111001100010;
mem[1299]=17'b11111111110000000;
mem[1300]=17'b00000000000010011;
mem[1301]=17'b11111000010010001;
mem[1302]=17'b00000000000001111;
mem[1303]=17'b11111001001111111;
mem[1304]=17'b11111110010110010;
mem[1305]=17'b00000000000000001;
mem[1306]=17'b00000000000000001;
mem[1307]=17'b11111100010000001;
mem[1308]=17'b00000000010110011;
mem[1309]=17'b11111111010111111;
mem[1310]=17'b00000000000000110;
mem[1311]=17'b00000001010110101;
mem[1312]=17'b11111110100001100;
mem[1313]=17'b00000010110011101;
mem[1314]=17'b11111110111001011;
mem[1315]=17'b01001101010111100;
mem[1316]=17'b00000000000001011;
mem[1317]=17'b11111100010011101;
mem[1318]=17'b11111111111010001;
mem[1319]=17'b00000000010000000;
mem[1320]=17'b00000000010011000;
mem[1321]=17'b11111111110110011;
mem[1322]=17'b11111110100111001;
mem[1323]=17'b00000000000011100;
mem[1324]=17'b00000000001100010;
mem[1325]=17'b11111111111100101;
mem[1326]=17'b00000000011011101;
mem[1327]=17'b00000001000111111;
mem[1328]=17'b11111110111111110;
mem[1329]=17'b11111110000011001;
mem[1330]=17'b00000000110101001;
mem[1331]=17'b00000001001111111;
mem[1332]=17'b11111110100101110;
mem[1333]=17'b11111111100101110;
mem[1334]=17'b11111111100001001;
mem[1335]=17'b11111111101101001;
mem[1336]=17'b11111110101111011;
mem[1337]=17'b00000000101100011;
mem[1338]=17'b11111011100011010;
mem[1339]=17'b11111001111000010;
mem[1340]=17'b00000010100111001;
mem[1341]=17'b11111111111000011;
mem[1342]=17'b11111111111010110;
mem[1343]=17'b11111101001111110;
mem[1344]=17'b11111001100010101;
mem[1345]=17'b00001010101101100;
mem[1346]=17'b00000001101000110;
mem[1347]=17'b00000000000010101;
mem[1348]=17'b11111111100000111;
mem[1349]=17'b00000000101010000;
mem[1350]=17'b00000000011110010;
mem[1351]=17'b11111111101101100;
mem[1352]=17'b00001011001001101;
mem[1353]=17'b00000000011111101;
mem[1354]=17'b11111111111011101;
mem[1355]=17'b00000000000110111;
mem[1356]=17'b00000000001001111;
mem[1357]=17'b11111111101011101;
mem[1358]=17'b11111111111110100;
mem[1359]=17'b00000000000100001;
mem[1360]=17'b00000000000011110;
mem[1361]=17'b00000000000001001;
mem[1362]=17'b00000000000000001;
mem[1363]=17'b00011011110111110;
mem[1364]=17'b00000000010101000;
mem[1365]=17'b00000000000110011;
mem[1366]=17'b11111111110010000;
mem[1367]=17'b00000000001000100;
mem[1368]=17'b00000000001011000;
mem[1369]=17'b11111111111100101;
mem[1370]=17'b00000000000000011;
mem[1371]=17'b11111110010011000;
mem[1372]=17'b00000000010101011;
mem[1373]=17'b11111110100100101;
mem[1374]=17'b11111100101111001;
mem[1375]=17'b00000000111101011;
mem[1376]=17'b11111110011111100;
mem[1377]=17'b11111101001000010;
mem[1378]=17'b00000000001011011;
mem[1379]=17'b11111111000111101;
mem[1380]=17'b11111111111101101;
mem[1381]=17'b11111111001111100;
mem[1382]=17'b00000000000001110;
mem[1383]=17'b11111111111111011;
mem[1384]=17'b11111001010010010;
mem[1385]=17'b11111111010010111;
mem[1386]=17'b00000001000000001;
mem[1387]=17'b00000011110000110;
mem[1388]=17'b11111111101110111;
mem[1389]=17'b00000000010110011;
mem[1390]=17'b11101100110111111;
mem[1391]=17'b11111011100011011;
mem[1392]=17'b11111100111000110;
mem[1393]=17'b00000001000100100;
mem[1394]=17'b11111011101001100;
mem[1395]=17'b11011110111000001;
mem[1396]=17'b00000000000010000;
mem[1397]=17'b11111110001110000;
mem[1398]=17'b00000000001011000;
mem[1399]=17'b11111111101110100;
mem[1400]=17'b11111111101110000;
mem[1401]=17'b11111111001101110;
mem[1402]=17'b11111001100110111;
mem[1403]=17'b11111111111111111;
mem[1404]=17'b00000000000110101;
mem[1405]=17'b11111111010100010;
mem[1406]=17'b00000000000010010;
mem[1407]=17'b00000000010100000;
mem[1408]=17'b11111110001110001;
mem[1409]=17'b00000000000101001;
mem[1410]=17'b00000001010110100;
mem[1411]=17'b00000000100101001;
mem[1412]=17'b00000000010001110;
mem[1413]=17'b11110000101001100;
mem[1414]=17'b11111111111101001;
mem[1415]=17'b11111110101111010;
mem[1416]=17'b11101001111111001;
mem[1417]=17'b00000000000011101;
mem[1418]=17'b00000000000000011;
mem[1419]=17'b11111011000001100;
mem[1420]=17'b00000110101000010;
mem[1421]=17'b00000000001010000;
mem[1422]=17'b00000000111100010;
mem[1423]=17'b00000000011110111;
mem[1424]=17'b00000000011000111;
mem[1425]=17'b00000000010000101;
mem[1426]=17'b00000000111001010;
mem[1427]=17'b11111111011110000;
mem[1428]=17'b00000000000001101;
mem[1429]=17'b11111100100100111;
mem[1430]=17'b11111111111100101;
mem[1431]=17'b11111011011010100;
mem[1432]=17'b00000000011101110;
mem[1433]=17'b00000011011000101;
mem[1434]=17'b11111110001101000;
mem[1435]=17'b11111101101000001;
mem[1436]=17'b00000000000010011;
mem[1437]=17'b00000001001011001;
mem[1438]=17'b11001110010100110;
mem[1439]=17'b00000010011100111;
mem[1440]=17'b00000000001010110;
mem[1441]=17'b00000000100000100;
mem[1442]=17'b11111101000010011;
mem[1443]=17'b11111110110101111;
mem[1444]=17'b00000000001001010;
mem[1445]=17'b11111100100011100;
mem[1446]=17'b00000001100100101;
mem[1447]=17'b11111111000011100;
mem[1448]=17'b00000000001010101;
mem[1449]=17'b00000001100010000;
mem[1450]=17'b11111111001011100;
mem[1451]=17'b00000000111110000;
mem[1452]=17'b00000000001100110;
mem[1453]=17'b11001001111101000;
mem[1454]=17'b11111101011000100;
mem[1455]=17'b11111110000111010;
mem[1456]=17'b11111111101100010;
mem[1457]=17'b00000001000100110;
mem[1458]=17'b00000000010100001;
mem[1459]=17'b00000000101111001;
mem[1460]=17'b00000001111000001;
mem[1461]=17'b00000010100011101;
mem[1462]=17'b11111111010101000;
mem[1463]=17'b00000000000101000;
mem[1464]=17'b00000000010011000;
mem[1465]=17'b11101110010000111;
mem[1466]=17'b11111111111111001;
mem[1467]=17'b11111111111111111;
mem[1468]=17'b00000001001011101;
mem[1469]=17'b00000000001110010;
mem[1470]=17'b00000000000001001;
mem[1471]=17'b00000000100000011;
mem[1472]=17'b00000010011111000;
mem[1473]=17'b00000101101010101;
mem[1474]=17'b00000001010100101;
mem[1475]=17'b00000001100111000;
mem[1476]=17'b11111111110001110;
mem[1477]=17'b00000010101001111;
mem[1478]=17'b00000000000110001;
mem[1479]=17'b00000010001111111;
mem[1480]=17'b11111111110100100;
mem[1481]=17'b00000001010101010;
mem[1482]=17'b00000101110010100;
mem[1483]=17'b11111011010100100;
mem[1484]=17'b11101110001011011;
mem[1485]=17'b11111101001100001;
mem[1486]=17'b00000001100111111;
mem[1487]=17'b11111111000000001;
mem[1488]=17'b00000000101000000;
mem[1489]=17'b00000001010110100;
mem[1490]=17'b11111111100001110;
mem[1491]=17'b11111110111011100;
mem[1492]=17'b11111100110011101;
mem[1493]=17'b00000000111101000;
mem[1494]=17'b11111111100000011;
mem[1495]=17'b11111111110111000;
mem[1496]=17'b11100011110001000;
mem[1497]=17'b00010101010011011;
mem[1498]=17'b11110101011100111;
mem[1499]=17'b11111111000011011;
mem[1500]=17'b00000000001100110;
mem[1501]=17'b00000001100110110;
mem[1502]=17'b00000000001011000;
mem[1503]=17'b00000000001011111;
mem[1504]=17'b11111111100000000;
mem[1505]=17'b11111111100100110;
mem[1506]=17'b11111111100100100;
mem[1507]=17'b11111110011110100;
mem[1508]=17'b00000000011100001;
mem[1509]=17'b00000000010000000;
mem[1510]=17'b11111110111110111;
mem[1511]=17'b11111111100000000;
mem[1512]=17'b11110000100010010;
mem[1513]=17'b11110111101101000;
mem[1514]=17'b00000000000001010;
mem[1515]=17'b00000000010000111;
mem[1516]=17'b11111110011000111;
mem[1517]=17'b00000011110011111;
mem[1518]=17'b11111000111111011;
mem[1519]=17'b00000001001001010;
mem[1520]=17'b11111101101011000;
mem[1521]=17'b00000000010010100;
mem[1522]=17'b11111111111100111;
mem[1523]=17'b11111111110101100;
mem[1524]=17'b00000000001101111;
mem[1525]=17'b00000000000010100;
mem[1526]=17'b00000000100101011;
mem[1527]=17'b00000101000100111;
mem[1528]=17'b11111111010111001;
mem[1529]=17'b00000001001010010;
mem[1530]=17'b11111110001100111;
mem[1531]=17'b11111111110001010;
mem[1532]=17'b11111111110001111;
mem[1533]=17'b00000000000001010;
mem[1534]=17'b11111110111110110;
mem[1535]=17'b00000000001010100;
mem[1536]=17'b00000001111111101;
mem[1537]=17'b11111000100001010;
mem[1538]=17'b00000000111110001;
mem[1539]=17'b11111111101000001;
mem[1540]=17'b00000011011000001;
mem[1541]=17'b11111110110101011;
mem[1542]=17'b11111111101101010;
mem[1543]=17'b11111111110001011;
mem[1544]=17'b11111111001001101;
mem[1545]=17'b11111110101001111;
mem[1546]=17'b00000010010001101;
mem[1547]=17'b00000001000010010;
mem[1548]=17'b11101000100000111;
mem[1549]=17'b00000101101111011;
mem[1550]=17'b00000000111101101;
mem[1551]=17'b00000000100010010;
mem[1552]=17'b00000001100111000;
mem[1553]=17'b00000000111101100;
mem[1554]=17'b11111111100011011;
mem[1555]=17'b11111101010000000;
mem[1556]=17'b11101011010100110;
mem[1557]=17'b11111110000111010;
mem[1558]=17'b00000000001010010;
mem[1559]=17'b11111111001010011;
mem[1560]=17'b00000010001100000;
mem[1561]=17'b11111111111000101;
mem[1562]=17'b11111111100101011;
mem[1563]=17'b00000000101001011;
mem[1564]=17'b00000000111110110;
mem[1565]=17'b11111001100010111;
mem[1566]=17'b11111110001101010;
mem[1567]=17'b00000011000100000;
mem[1568]=17'b00000000011010101;
mem[1569]=17'b00000001000000110;
mem[1570]=17'b11111111010000100;
mem[1571]=17'b11111101100100010;
mem[1572]=17'b00000000111011001;
mem[1573]=17'b11111111111101011;
mem[1574]=17'b11111101000100101;
mem[1575]=17'b00000000101010011;
mem[1576]=17'b00000000101111101;
mem[1577]=17'b00000000001010100;
mem[1578]=17'b11111101101110000;
mem[1579]=17'b11111111000110000;
mem[1580]=17'b00000001000001101;
mem[1581]=17'b00000001111110001;
mem[1582]=17'b00000111011001011;
mem[1583]=17'b00000000111011100;
mem[1584]=17'b11111111001001100;
mem[1585]=17'b11111111111001111;
mem[1586]=17'b00000000101111001;
mem[1587]=17'b11111101111111010;
mem[1588]=17'b11111111111100001;
mem[1589]=17'b11111111101101100;
mem[1590]=17'b00000000010101001;
mem[1591]=17'b11111110011011101;
mem[1592]=17'b11111110111110100;
mem[1593]=17'b11111000100111111;
mem[1594]=17'b00000000000011000;
mem[1595]=17'b11111111111111111;
mem[1596]=17'b00000000011100010;
mem[1597]=17'b11111111110001010;
mem[1598]=17'b00000000111111111;
mem[1599]=17'b11111111101101010;
mem[1600]=17'b11111111110000110;
mem[1601]=17'b11111111000110100;
mem[1602]=17'b00000000000001111;
mem[1603]=17'b00000000100001110;
mem[1604]=17'b11111111111100010;
mem[1605]=17'b00000000010010001;
mem[1606]=17'b00001111111000101;
mem[1607]=17'b00001111111111001;
mem[1608]=17'b00000010001101111;
mem[1609]=17'b00000000000010000;
mem[1610]=17'b11111110111011110;
mem[1611]=17'b00000000001110011;
mem[1612]=17'b11111011100110111;
mem[1613]=17'b11111111111101010;
mem[1614]=17'b00000000000010100;
mem[1615]=17'b11111011101001111;
mem[1616]=17'b11111111110101010;
mem[1617]=17'b11111111111010100;
mem[1618]=17'b00000000010011010;
mem[1619]=17'b11111111010010100;
mem[1620]=17'b00000000000110001;
mem[1621]=17'b11111110110010111;
mem[1622]=17'b11111101101010110;
mem[1623]=17'b11111111011011010;
mem[1624]=17'b00000011011010010;
mem[1625]=17'b11111101010101001;
mem[1626]=17'b11111111111011000;
mem[1627]=17'b00000000100111000;
mem[1628]=17'b11111111001000010;
mem[1629]=17'b00000001001000100;
mem[1630]=17'b00000000000000110;
mem[1631]=17'b00000111010110001;
mem[1632]=17'b00000001101110110;
mem[1633]=17'b11100001010000100;
mem[1634]=17'b11111111111010110;
mem[1635]=17'b11111111101111111;
mem[1636]=17'b11111111010010101;
mem[1637]=17'b00000000000000011;
mem[1638]=17'b00000000010000110;
mem[1639]=17'b11111111101111000;
mem[1640]=17'b00000100001011001;
mem[1641]=17'b11111110011111011;
mem[1642]=17'b00000100110101100;
mem[1643]=17'b11111111011010100;
mem[1644]=17'b00001011100000101;
mem[1645]=17'b11111111110001100;
mem[1646]=17'b00000011010111010;
mem[1647]=17'b00000001000000101;
mem[1648]=17'b11111111000101011;
mem[1649]=17'b00000000010101100;
mem[1650]=17'b11111111101010111;
mem[1651]=17'b11111100001000001;
mem[1652]=17'b00000010000100110;
mem[1653]=17'b00000000000001111;
mem[1654]=17'b11110111011001111;
mem[1655]=17'b00000001101010010;
mem[1656]=17'b11111111001011010;
mem[1657]=17'b00000000010110010;
mem[1658]=17'b00000000000001100;
mem[1659]=17'b00000000000010011;
mem[1660]=17'b00000001000111001;
mem[1661]=17'b11111110011001111;
mem[1662]=17'b00000000000111110;
mem[1663]=17'b11111111111101001;
mem[1664]=17'b00000000000101100;
mem[1665]=17'b00000000000011110;
mem[1666]=17'b00000010000100000;
mem[1667]=17'b11111110011101010;
mem[1668]=17'b11111111000100001;
mem[1669]=17'b11111110111111001;
mem[1670]=17'b00000000011100110;
mem[1671]=17'b00000000001010101;
mem[1672]=17'b11110111101111101;
mem[1673]=17'b11111111111001100;
mem[1674]=17'b00000000010000000;
mem[1675]=17'b00000001100110011;
mem[1676]=17'b11111111110000111;
mem[1677]=17'b00000000000111111;
mem[1678]=17'b00000001010101100;
mem[1679]=17'b11111111010000101;
mem[1680]=17'b11111000000011011;
mem[1681]=17'b00000000010010000;
mem[1682]=17'b00000000000101000;
mem[1683]=17'b11111111100111110;
mem[1684]=17'b11111101001101010;
mem[1685]=17'b11101011110011001;
mem[1686]=17'b11111100100010000;
mem[1687]=17'b00000000000001111;
mem[1688]=17'b00011010111000001;
mem[1689]=17'b11111011000101011;
mem[1690]=17'b11111111001110110;
mem[1691]=17'b11111111100010011;
mem[1692]=17'b11111111000010000;
mem[1693]=17'b00000000011111100;
mem[1694]=17'b00001001000110010;
mem[1695]=17'b11111011111100000;
mem[1696]=17'b00000000000011011;
mem[1697]=17'b11111111101000110;
mem[1698]=17'b11111110101111011;
mem[1699]=17'b11111111111101000;
mem[1700]=17'b11111111110010111;
mem[1701]=17'b00000000000010010;
mem[1702]=17'b11110011101110000;
mem[1703]=17'b11110010000101111;
mem[1704]=17'b11110001111001001;
mem[1705]=17'b00000000011111010;
mem[1706]=17'b00000000010011110;
mem[1707]=17'b11111011001110000;
mem[1708]=17'b11111101100000101;
mem[1709]=17'b11111111111101011;
mem[1710]=17'b00000000000000011;
mem[1711]=17'b00000010010110101;
mem[1712]=17'b00000101011010000;
mem[1713]=17'b11111111111111101;
mem[1714]=17'b00000000011001100;
mem[1715]=17'b00000000111001111;
mem[1716]=17'b00000000000110001;
mem[1717]=17'b00000000001111000;
mem[1718]=17'b00000000001100001;
mem[1719]=17'b00000000000000001;
mem[1720]=17'b11111111111000010;
mem[1721]=17'b00000000101010100;
mem[1722]=17'b11111111110001111;
mem[1723]=17'b11111111101101110;
mem[1724]=17'b00000000011010100;
mem[1725]=17'b11111111111110000;
mem[1726]=17'b00000001110001000;
mem[1727]=17'b11111101111001000;
mem[1728]=17'b11111111100011000;
mem[1729]=17'b11111111110101010;
mem[1730]=17'b00000000001111011;
mem[1731]=17'b00000000100001111;
mem[1732]=17'b11111111110010000;
mem[1733]=17'b00000000000110010;
mem[1734]=17'b11110111001110001;
mem[1735]=17'b00000110111100000;
mem[1736]=17'b11111111011100111;
mem[1737]=17'b00000000101010101;
mem[1738]=17'b11111011111111100;
mem[1739]=17'b00000000010001010;
mem[1740]=17'b00000000100110000;
mem[1741]=17'b00000001010000101;
mem[1742]=17'b11111101011010100;
mem[1743]=17'b00000000110011011;
mem[1744]=17'b11111111011110010;
mem[1745]=17'b00000010110010001;
mem[1746]=17'b11111111111010010;
mem[1747]=17'b00000000000011001;
mem[1748]=17'b00000000011101000;
mem[1749]=17'b00000000011110110;
mem[1750]=17'b11111111111111101;
mem[1751]=17'b11111110100000001;
mem[1752]=17'b11111100011111111;
mem[1753]=17'b00011100100100000;
mem[1754]=17'b00000001000110110;
mem[1755]=17'b11111111110011110;
mem[1756]=17'b11111111100110000;
mem[1757]=17'b00000000010101010;
mem[1758]=17'b11111111011000001;
mem[1759]=17'b11111110101110001;
mem[1760]=17'b00000000000100000;
mem[1761]=17'b11111100010110111;
mem[1762]=17'b00000001110000100;
mem[1763]=17'b11111111001001110;
mem[1764]=17'b00000001111100010;
mem[1765]=17'b11111111001101000;
mem[1766]=17'b11111100101001010;
mem[1767]=17'b00000011101001111;
mem[1768]=17'b00000001001000110;
mem[1769]=17'b11111111110010011;
mem[1770]=17'b11111111010000101;
mem[1771]=17'b11111111111101011;
mem[1772]=17'b00000000001101101;
mem[1773]=17'b00000000101110000;
mem[1774]=17'b11111110111101110;
mem[1775]=17'b11111111111100110;
mem[1776]=17'b00000001010001010;
mem[1777]=17'b11111111111010011;
mem[1778]=17'b00000000001001100;
mem[1779]=17'b11111111010011001;
mem[1780]=17'b11111101011111100;
mem[1781]=17'b00000001111001100;
mem[1782]=17'b00000010100101111;
mem[1783]=17'b00000000111100011;
mem[1784]=17'b11111111100010100;
mem[1785]=17'b11111111011011111;
mem[1786]=17'b11111111101101110;
mem[1787]=17'b00000000011000110;
mem[1788]=17'b00000000000011010;
mem[1789]=17'b00000000001010000;
mem[1790]=17'b11111100000101111;
mem[1791]=17'b00000000000101100;
mem[1792]=17'b00000100010010100;
mem[1793]=17'b00000000000111100;
mem[1794]=17'b11111010110001010;
mem[1795]=17'b11111101001101011;
mem[1796]=17'b11111110101110100;
mem[1797]=17'b11111110010010100;
mem[1798]=17'b00000000001100010;
mem[1799]=17'b00000000001001110;
mem[1800]=17'b11111110010111011;
mem[1801]=17'b11111110000111110;
mem[1802]=17'b00000000111101011;
mem[1803]=17'b11111111010010011;
mem[1804]=17'b00000000110100001;
mem[1805]=17'b00000000010000000;
mem[1806]=17'b11111111011010111;
mem[1807]=17'b11111111100000111;
mem[1808]=17'b00000100111101110;
mem[1809]=17'b11110110001110110;
mem[1810]=17'b11111111101011100;
mem[1811]=17'b11101100100110011;
mem[1812]=17'b00000000001110010;
mem[1813]=17'b11111111101111011;
mem[1814]=17'b00000000000101110;
mem[1815]=17'b11111111111000000;
mem[1816]=17'b00000000000001110;
mem[1817]=17'b11111100101101010;
mem[1818]=17'b00000010101011001;
mem[1819]=17'b00000000000001010;
mem[1820]=17'b11111110111001010;
mem[1821]=17'b11111111011110100;
mem[1822]=17'b00000001000001000;
mem[1823]=17'b00001111111101101;
mem[1824]=17'b11101100001010000;
mem[1825]=17'b11111111110111110;
mem[1826]=17'b11111100001100111;
mem[1827]=17'b00000011011110000;
mem[1828]=17'b00000000000111000;
mem[1829]=17'b00000000011001101;
mem[1830]=17'b11111110011100101;
mem[1831]=17'b00001010001011001;
mem[1832]=17'b11111111100010110;
mem[1833]=17'b11111111111110000;
mem[1834]=17'b00010101000010011;
mem[1835]=17'b00000000100010110;
mem[1836]=17'b00001001101010101;
mem[1837]=17'b00000000001100010;
mem[1838]=17'b11111010111011010;
mem[1839]=17'b00001010011111011;
mem[1840]=17'b11111101100001110;
mem[1841]=17'b11100010110100101;
mem[1842]=17'b11111100110100011;
mem[1843]=17'b00000000000101000;
mem[1844]=17'b11111110111100111;
mem[1845]=17'b11111110111111100;
mem[1846]=17'b00000000100110001;
mem[1847]=17'b11111110100010110;
mem[1848]=17'b00000000010011010;
mem[1849]=17'b11111110001000101;
mem[1850]=17'b00000101101110111;
mem[1851]=17'b00100010000010100;
mem[1852]=17'b11111111010110011;
mem[1853]=17'b00000000000111001;
mem[1854]=17'b01001000100001000;
mem[1855]=17'b11111101101011011;
mem[1856]=17'b11111111001011111;
mem[1857]=17'b00000000000111010;
mem[1858]=17'b00000000001000101;
mem[1859]=17'b00000000001000000;
mem[1860]=17'b00000000001111111;
mem[1861]=17'b11111111000011011;
mem[1862]=17'b11111110101101010;
mem[1863]=17'b00000000000100011;
mem[1864]=17'b00000000000010000;
mem[1865]=17'b00000001111111101;
mem[1866]=17'b11111111111010110;
mem[1867]=17'b11111111111011100;
mem[1868]=17'b00000000000101001;
mem[1869]=17'b11111111110101100;
mem[1870]=17'b00000001001100000;
mem[1871]=17'b11111011101001101;
mem[1872]=17'b11111101000110000;
mem[1873]=17'b11110111111001100;
mem[1874]=17'b11111111111000101;
mem[1875]=17'b00000001000110100;
mem[1876]=17'b11111110110010100;
mem[1877]=17'b00010010111010000;
mem[1878]=17'b00000000111100100;
mem[1879]=17'b11111111111001011;
mem[1880]=17'b11111111011111100;
mem[1881]=17'b11111010110010010;
mem[1882]=17'b11111110111010000;
mem[1883]=17'b00000001000001101;
mem[1884]=17'b00000000000110001;
mem[1885]=17'b11111111100101000;
mem[1886]=17'b11111101010111011;
mem[1887]=17'b11111111000010101;
mem[1888]=17'b00000001010110011;
mem[1889]=17'b00000000010010101;
mem[1890]=17'b00000000111100111;
mem[1891]=17'b00000001010111001;
mem[1892]=17'b00000000101110110;
mem[1893]=17'b00000100010010100;
mem[1894]=17'b00000000110101010;
mem[1895]=17'b00000001101110101;
mem[1896]=17'b11111111111011100;
mem[1897]=17'b00000000001101110;
mem[1898]=17'b00000001001001111;
mem[1899]=17'b00000000010100000;
mem[1900]=17'b11111111100111011;
mem[1901]=17'b11111110011011000;
mem[1902]=17'b11111111100011101;
mem[1903]=17'b00000000011000010;
mem[1904]=17'b00000000100011010;
mem[1905]=17'b00000001000010010;
mem[1906]=17'b11111111110100100;
mem[1907]=17'b00000001000010010;
mem[1908]=17'b11111101111110101;
mem[1909]=17'b11111100010001110;
mem[1910]=17'b00000001001011110;
mem[1911]=17'b11111110101111100;
mem[1912]=17'b00000001010011101;
mem[1913]=17'b00000000001101111;
mem[1914]=17'b11111011011111100;
mem[1915]=17'b11111111011001101;
mem[1916]=17'b00000001011111101;
mem[1917]=17'b00000101001110111;
mem[1918]=17'b00000000001100000;
mem[1919]=17'b00000110101011000;
mem[1920]=17'b11111100111110100;
mem[1921]=17'b00000000001100101;
mem[1922]=17'b11101100111110001;
mem[1923]=17'b00000001010000010;
mem[1924]=17'b00000000000011110;
mem[1925]=17'b00000000001111000;
mem[1926]=17'b00000000000000100;
mem[1927]=17'b11111111111111101;
mem[1928]=17'b00000000100110011;
mem[1929]=17'b11111101111001100;
mem[1930]=17'b00000001101010110;
mem[1931]=17'b11111111010111110;
mem[1932]=17'b11111111111111111;
mem[1933]=17'b11111111111010101;
mem[1934]=17'b00000000000001111;
mem[1935]=17'b00001110010011111;
mem[1936]=17'b00000000001010110;
mem[1937]=17'b00001100100110001;
mem[1938]=17'b11111111010100110;
mem[1939]=17'b11111111111110100;
mem[1940]=17'b11111111111001001;
mem[1941]=17'b11111111101000100;
mem[1942]=17'b11111111111010100;
mem[1943]=17'b11111111100001011;
mem[1944]=17'b11101100001111100;
mem[1945]=17'b00000000101000101;
mem[1946]=17'b00000000000100001;
mem[1947]=17'b11111001011111100;
mem[1948]=17'b11111110011100110;
mem[1949]=17'b00000011001101001;
mem[1950]=17'b00000000000000000;
mem[1951]=17'b00000001011101111;
mem[1952]=17'b11111111101010011;
mem[1953]=17'b00000000011110110;
mem[1954]=17'b11111110111001010;
mem[1955]=17'b11111111011110001;
mem[1956]=17'b00000010010000100;
mem[1957]=17'b11111111110111100;
mem[1958]=17'b00000000010010011;
mem[1959]=17'b00000000011111100;
mem[1960]=17'b00000000000100001;
mem[1961]=17'b11111001010010100;
mem[1962]=17'b00000011101101010;
mem[1963]=17'b11111111111100010;
mem[1964]=17'b11111111111010010;
mem[1965]=17'b11111101111110000;
mem[1966]=17'b11111111111111110;
mem[1967]=17'b00000000000000111;
mem[1968]=17'b11111110100111011;
mem[1969]=17'b11111110011101100;
mem[1970]=17'b11111110100010100;
mem[1971]=17'b00000000011001001;
mem[1972]=17'b00000001011011101;
mem[1973]=17'b11111011001011111;
mem[1974]=17'b11111011110010111;
mem[1975]=17'b00000000000100100;
mem[1976]=17'b11111100100011101;
mem[1977]=17'b11111110011011011;
mem[1978]=17'b11111111111010011;
mem[1979]=17'b00000001000111000;
mem[1980]=17'b11111110100111001;
mem[1981]=17'b00000000000001101;
mem[1982]=17'b11110110110100110;
mem[1983]=17'b11111011101011110;
mem[1984]=17'b11111011111101011;
mem[1985]=17'b00000001001010111;
mem[1986]=17'b11111111111111011;
mem[1987]=17'b11111111110001011;
mem[1988]=17'b00000000011001011;
mem[1989]=17'b11111110111100101;
mem[1990]=17'b00000000010000001;
mem[1991]=17'b11111110101111100;
mem[1992]=17'b00000000001000100;
mem[1993]=17'b11111111110010101;
mem[1994]=17'b11111111111010011;
mem[1995]=17'b00000000001111000;
mem[1996]=17'b00000001000011001;
mem[1997]=17'b11111011000110000;
mem[1998]=17'b00000000001001011;
mem[1999]=17'b00000000010010001;
mem[2000]=17'b11111111100001001;
mem[2001]=17'b11111111110000100;
mem[2002]=17'b11111111110000001;
mem[2003]=17'b00000001001111010;
mem[2004]=17'b11111111101010110;
mem[2005]=17'b11111010100010011;
mem[2006]=17'b11111111101011110;
mem[2007]=17'b11111111101100010;
mem[2008]=17'b00000000000100111;
mem[2009]=17'b11111101000100010;
mem[2010]=17'b00000001101000011;
mem[2011]=17'b00000000001110001;
mem[2012]=17'b11111110100011001;
mem[2013]=17'b11111111111101000;
mem[2014]=17'b11111111111101001;
mem[2015]=17'b00000001000111010;
mem[2016]=17'b00000110000111111;
mem[2017]=17'b00000000001011110;
mem[2018]=17'b11111111111111100;
mem[2019]=17'b11111110101011000;
mem[2020]=17'b00001000101001001;
mem[2021]=17'b00000000011100100;
mem[2022]=17'b00000000101000101;
mem[2023]=17'b11111111111101110;
mem[2024]=17'b11111110111100010;
mem[2025]=17'b00000000010000010;
mem[2026]=17'b00000000110111100;
mem[2027]=17'b00000001101101000;
mem[2028]=17'b11111111110100000;
mem[2029]=17'b00000000010001011;
mem[2030]=17'b00000000000101101;
mem[2031]=17'b00000000010001000;
mem[2032]=17'b11111111111000010;
mem[2033]=17'b11111111100001110;
mem[2034]=17'b00000000001101101;
mem[2035]=17'b00000000011100000;
mem[2036]=17'b00000001000110010;
mem[2037]=17'b11110000111011011;
mem[2038]=17'b00000101000001101;
mem[2039]=17'b11111111111111101;
mem[2040]=17'b11111111111000101;
mem[2041]=17'b11111111011110000;
mem[2042]=17'b11111111101110011;
mem[2043]=17'b00000000001111110;
mem[2044]=17'b11111111111111111;
mem[2045]=17'b11111101011100000;
mem[2046]=17'b00000100100100100;
mem[2047]=17'b00000000001010100;
mem[2048]=17'b00000010100011011;
mem[2049]=17'b11110101111111011;
mem[2050]=17'b00000011001001111;
mem[2051]=17'b11111100010011010;
mem[2052]=17'b00000000011111100;
mem[2053]=17'b00001100100101010;
mem[2054]=17'b11111111111111110;
mem[2055]=17'b00000000011011000;
mem[2056]=17'b11111100101011001;
mem[2057]=17'b11111111011011001;
mem[2058]=17'b00001111010110110;
mem[2059]=17'b00000000110010001;
mem[2060]=17'b11110001011101111;
mem[2061]=17'b01101100000101000;
mem[2062]=17'b00000000100101110;
mem[2063]=17'b00000000101100001;
mem[2064]=17'b11111111111010101;
mem[2065]=17'b00000000101010010;
mem[2066]=17'b00000000000110000;
mem[2067]=17'b11111010110100001;
mem[2068]=17'b11111111011010000;
mem[2069]=17'b00000001001010111;
mem[2070]=17'b11110110110011101;
mem[2071]=17'b00011111001011000;
mem[2072]=17'b00000011000010000;
mem[2073]=17'b11111111110010100;
mem[2074]=17'b00000001010101000;
mem[2075]=17'b11111101100011100;
mem[2076]=17'b00000001001000010;
mem[2077]=17'b00000000010000100;
mem[2078]=17'b00000010001010000;
mem[2079]=17'b00000000100100101;
mem[2080]=17'b00000000100100101;
mem[2081]=17'b11111110111101100;
mem[2082]=17'b00000001000100110;
mem[2083]=17'b11111101000100101;
mem[2084]=17'b11111111111111111;
mem[2085]=17'b11111111111110100;
mem[2086]=17'b00000011011001100;
mem[2087]=17'b11111000111110111;
mem[2088]=17'b00000000011110111;
mem[2089]=17'b11111111110011110;
mem[2090]=17'b00000000000010000;
mem[2091]=17'b11111011110001100;
mem[2092]=17'b00000000001011001;
mem[2093]=17'b11111010011010011;
mem[2094]=17'b00000001010110001;
mem[2095]=17'b00000100101001111;
mem[2096]=17'b11111101101011000;
mem[2097]=17'b00000011001001110;
mem[2098]=17'b11111111101110101;
mem[2099]=17'b11111111110101101;
mem[2100]=17'b11111111111000011;
mem[2101]=17'b00000000000110010;
mem[2102]=17'b00000000011110000;
mem[2103]=17'b11111110001101110;
mem[2104]=17'b11111101001101111;
mem[2105]=17'b00000000001101000;
mem[2106]=17'b11111111011100111;
mem[2107]=17'b11111100110000110;
mem[2108]=17'b00000000110111011;
mem[2109]=17'b00000000000111011;
mem[2110]=17'b11111111100011010;
mem[2111]=17'b00000000011101101;
mem[2112]=17'b00000001110000001;
mem[2113]=17'b11111111111101010;
mem[2114]=17'b11111110100000111;
mem[2115]=17'b11111111100010011;
mem[2116]=17'b11111111100101001;
mem[2117]=17'b00000000000101111;
mem[2118]=17'b00000000001101100;
mem[2119]=17'b00000000001011001;
mem[2120]=17'b00000000000100010;
mem[2121]=17'b11111111101101000;
mem[2122]=17'b00000000100110101;
mem[2123]=17'b00000001000000010;
mem[2124]=17'b11111111111000101;
mem[2125]=17'b00001001000001110;
mem[2126]=17'b11111111110010010;
mem[2127]=17'b00000000000010000;
mem[2128]=17'b11111100001000010;
mem[2129]=17'b00101001011100110;
mem[2130]=17'b11111111111010110;
mem[2131]=17'b00000000011100111;
mem[2132]=17'b11111110101001010;
mem[2133]=17'b00000010001110110;
mem[2134]=17'b00001000101000011;
end

always@(posedge clk)
begin
  if (we) begin
    mem[addr] <= din;
  end
end

always @(posedge clk) dout <= mem[addr];

endmodule
